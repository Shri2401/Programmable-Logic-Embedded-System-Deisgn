`timescale 1 ns/100 ps
// Version: v12.6 12.900.20.24


module MSS_010(
       CAN_RXBUS_MGPIO3A_H2F_A,
       CAN_RXBUS_MGPIO3A_H2F_B,
       CAN_TX_EBL_MGPIO4A_H2F_A,
       CAN_TX_EBL_MGPIO4A_H2F_B,
       CAN_TXBUS_MGPIO2A_H2F_A,
       CAN_TXBUS_MGPIO2A_H2F_B,
       CLK_CONFIG_APB,
       COMMS_INT,
       CONFIG_PRESET_N,
       EDAC_ERROR,
       F_FM0_RDATA,
       F_FM0_READYOUT,
       F_FM0_RESP,
       F_HM0_ADDR,
       F_HM0_ENABLE,
       F_HM0_SEL,
       F_HM0_SIZE,
       F_HM0_TRANS1,
       F_HM0_WDATA,
       F_HM0_WRITE,
       FAB_CHRGVBUS,
       FAB_DISCHRGVBUS,
       FAB_DMPULLDOWN,
       FAB_DPPULLDOWN,
       FAB_DRVVBUS,
       FAB_IDPULLUP,
       FAB_OPMODE,
       FAB_SUSPENDM,
       FAB_TERMSEL,
       FAB_TXVALID,
       FAB_VCONTROL,
       FAB_VCONTROLLOADM,
       FAB_XCVRSEL,
       FAB_XDATAOUT,
       FACC_GLMUX_SEL,
       FIC32_0_MASTER,
       FIC32_1_MASTER,
       FPGA_RESET_N,
       GTX_CLK,
       H2F_INTERRUPT,
       H2F_NMI,
       H2FCALIB,
       I2C0_SCL_MGPIO31B_H2F_A,
       I2C0_SCL_MGPIO31B_H2F_B,
       I2C0_SDA_MGPIO30B_H2F_A,
       I2C0_SDA_MGPIO30B_H2F_B,
       I2C1_SCL_MGPIO1A_H2F_A,
       I2C1_SCL_MGPIO1A_H2F_B,
       I2C1_SDA_MGPIO0A_H2F_A,
       I2C1_SDA_MGPIO0A_H2F_B,
       MDCF,
       MDOENF,
       MDOF,
       MMUART0_CTS_MGPIO19B_H2F_A,
       MMUART0_CTS_MGPIO19B_H2F_B,
       MMUART0_DCD_MGPIO22B_H2F_A,
       MMUART0_DCD_MGPIO22B_H2F_B,
       MMUART0_DSR_MGPIO20B_H2F_A,
       MMUART0_DSR_MGPIO20B_H2F_B,
       MMUART0_DTR_MGPIO18B_H2F_A,
       MMUART0_DTR_MGPIO18B_H2F_B,
       MMUART0_RI_MGPIO21B_H2F_A,
       MMUART0_RI_MGPIO21B_H2F_B,
       MMUART0_RTS_MGPIO17B_H2F_A,
       MMUART0_RTS_MGPIO17B_H2F_B,
       MMUART0_RXD_MGPIO28B_H2F_A,
       MMUART0_RXD_MGPIO28B_H2F_B,
       MMUART0_SCK_MGPIO29B_H2F_A,
       MMUART0_SCK_MGPIO29B_H2F_B,
       MMUART0_TXD_MGPIO27B_H2F_A,
       MMUART0_TXD_MGPIO27B_H2F_B,
       MMUART1_DTR_MGPIO12B_H2F_A,
       MMUART1_RTS_MGPIO11B_H2F_A,
       MMUART1_RTS_MGPIO11B_H2F_B,
       MMUART1_RXD_MGPIO26B_H2F_A,
       MMUART1_RXD_MGPIO26B_H2F_B,
       MMUART1_SCK_MGPIO25B_H2F_A,
       MMUART1_SCK_MGPIO25B_H2F_B,
       MMUART1_TXD_MGPIO24B_H2F_A,
       MMUART1_TXD_MGPIO24B_H2F_B,
       MPLL_LOCK,
       PER2_FABRIC_PADDR,
       PER2_FABRIC_PENABLE,
       PER2_FABRIC_PSEL,
       PER2_FABRIC_PWDATA,
       PER2_FABRIC_PWRITE,
       RTC_MATCH,
       SLEEPDEEP,
       SLEEPHOLDACK,
       SLEEPING,
       SMBALERT_NO0,
       SMBALERT_NO1,
       SMBSUS_NO0,
       SMBSUS_NO1,
       SPI0_CLK_OUT,
       SPI0_SDI_MGPIO5A_H2F_A,
       SPI0_SDI_MGPIO5A_H2F_B,
       SPI0_SDO_MGPIO6A_H2F_A,
       SPI0_SDO_MGPIO6A_H2F_B,
       SPI0_SS0_MGPIO7A_H2F_A,
       SPI0_SS0_MGPIO7A_H2F_B,
       SPI0_SS1_MGPIO8A_H2F_A,
       SPI0_SS1_MGPIO8A_H2F_B,
       SPI0_SS2_MGPIO9A_H2F_A,
       SPI0_SS2_MGPIO9A_H2F_B,
       SPI0_SS3_MGPIO10A_H2F_A,
       SPI0_SS3_MGPIO10A_H2F_B,
       SPI0_SS4_MGPIO19A_H2F_A,
       SPI0_SS5_MGPIO20A_H2F_A,
       SPI0_SS6_MGPIO21A_H2F_A,
       SPI0_SS7_MGPIO22A_H2F_A,
       SPI1_CLK_OUT,
       SPI1_SDI_MGPIO11A_H2F_A,
       SPI1_SDI_MGPIO11A_H2F_B,
       SPI1_SDO_MGPIO12A_H2F_A,
       SPI1_SDO_MGPIO12A_H2F_B,
       SPI1_SS0_MGPIO13A_H2F_A,
       SPI1_SS0_MGPIO13A_H2F_B,
       SPI1_SS1_MGPIO14A_H2F_A,
       SPI1_SS1_MGPIO14A_H2F_B,
       SPI1_SS2_MGPIO15A_H2F_A,
       SPI1_SS2_MGPIO15A_H2F_B,
       SPI1_SS3_MGPIO16A_H2F_A,
       SPI1_SS3_MGPIO16A_H2F_B,
       SPI1_SS4_MGPIO17A_H2F_A,
       SPI1_SS5_MGPIO18A_H2F_A,
       SPI1_SS6_MGPIO23A_H2F_A,
       SPI1_SS7_MGPIO24A_H2F_A,
       TCGF,
       TRACECLK,
       TRACEDATA,
       TX_CLK,
       TX_ENF,
       TX_ERRF,
       TXCTL_EN_RIF,
       TXD_RIF,
       TXDF,
       TXEV,
       WDOGTIMEOUT,
       F_ARREADY_HREADYOUT1,
       F_AWREADY_HREADYOUT0,
       F_BID,
       F_BRESP_HRESP0,
       F_BVALID,
       F_RDATA_HRDATA01,
       F_RID,
       F_RLAST,
       F_RRESP_HRESP1,
       F_RVALID,
       F_WREADY,
       MDDR_FABRIC_PRDATA,
       MDDR_FABRIC_PREADY,
       MDDR_FABRIC_PSLVERR,
       CAN_RXBUS_F2H_SCP,
       CAN_TX_EBL_F2H_SCP,
       CAN_TXBUS_F2H_SCP,
       COLF,
       CRSF,
       F2_DMAREADY,
       F2H_INTERRUPT,
       F2HCALIB,
       F_DMAREADY,
       F_FM0_ADDR,
       F_FM0_ENABLE,
       F_FM0_MASTLOCK,
       F_FM0_READY,
       F_FM0_SEL,
       F_FM0_SIZE,
       F_FM0_TRANS1,
       F_FM0_WDATA,
       F_FM0_WRITE,
       F_HM0_RDATA,
       F_HM0_READY,
       F_HM0_RESP,
       FAB_AVALID,
       FAB_HOSTDISCON,
       FAB_IDDIG,
       FAB_LINESTATE,
       FAB_M3_RESET_N,
       FAB_PLL_LOCK,
       FAB_RXACTIVE,
       FAB_RXERROR,
       FAB_RXVALID,
       FAB_RXVALIDH,
       FAB_SESSEND,
       FAB_TXREADY,
       FAB_VBUSVALID,
       FAB_VSTATUS,
       FAB_XDATAIN,
       GTX_CLKPF,
       I2C0_BCLK,
       I2C0_SCL_F2H_SCP,
       I2C0_SDA_F2H_SCP,
       I2C1_BCLK,
       I2C1_SCL_F2H_SCP,
       I2C1_SDA_F2H_SCP,
       MDIF,
       MGPIO0A_F2H_GPIN,
       MGPIO10A_F2H_GPIN,
       MGPIO11A_F2H_GPIN,
       MGPIO11B_F2H_GPIN,
       MGPIO12A_F2H_GPIN,
       MGPIO13A_F2H_GPIN,
       MGPIO14A_F2H_GPIN,
       MGPIO15A_F2H_GPIN,
       MGPIO16A_F2H_GPIN,
       MGPIO17B_F2H_GPIN,
       MGPIO18B_F2H_GPIN,
       MGPIO19B_F2H_GPIN,
       MGPIO1A_F2H_GPIN,
       MGPIO20B_F2H_GPIN,
       MGPIO21B_F2H_GPIN,
       MGPIO22B_F2H_GPIN,
       MGPIO24B_F2H_GPIN,
       MGPIO25B_F2H_GPIN,
       MGPIO26B_F2H_GPIN,
       MGPIO27B_F2H_GPIN,
       MGPIO28B_F2H_GPIN,
       MGPIO29B_F2H_GPIN,
       MGPIO2A_F2H_GPIN,
       MGPIO30B_F2H_GPIN,
       MGPIO31B_F2H_GPIN,
       MGPIO3A_F2H_GPIN,
       MGPIO4A_F2H_GPIN,
       MGPIO5A_F2H_GPIN,
       MGPIO6A_F2H_GPIN,
       MGPIO7A_F2H_GPIN,
       MGPIO8A_F2H_GPIN,
       MGPIO9A_F2H_GPIN,
       MMUART0_CTS_F2H_SCP,
       MMUART0_DCD_F2H_SCP,
       MMUART0_DSR_F2H_SCP,
       MMUART0_DTR_F2H_SCP,
       MMUART0_RI_F2H_SCP,
       MMUART0_RTS_F2H_SCP,
       MMUART0_RXD_F2H_SCP,
       MMUART0_SCK_F2H_SCP,
       MMUART0_TXD_F2H_SCP,
       MMUART1_CTS_F2H_SCP,
       MMUART1_DCD_F2H_SCP,
       MMUART1_DSR_F2H_SCP,
       MMUART1_RI_F2H_SCP,
       MMUART1_RTS_F2H_SCP,
       MMUART1_RXD_F2H_SCP,
       MMUART1_SCK_F2H_SCP,
       MMUART1_TXD_F2H_SCP,
       PER2_FABRIC_PRDATA,
       PER2_FABRIC_PREADY,
       PER2_FABRIC_PSLVERR,
       RCGF,
       RX_CLKPF,
       RX_DVF,
       RX_ERRF,
       RX_EV,
       RXDF,
       SLEEPHOLDREQ,
       SMBALERT_NI0,
       SMBALERT_NI1,
       SMBSUS_NI0,
       SMBSUS_NI1,
       SPI0_CLK_IN,
       SPI0_SDI_F2H_SCP,
       SPI0_SDO_F2H_SCP,
       SPI0_SS0_F2H_SCP,
       SPI0_SS1_F2H_SCP,
       SPI0_SS2_F2H_SCP,
       SPI0_SS3_F2H_SCP,
       SPI1_CLK_IN,
       SPI1_SDI_F2H_SCP,
       SPI1_SDO_F2H_SCP,
       SPI1_SS0_F2H_SCP,
       SPI1_SS1_F2H_SCP,
       SPI1_SS2_F2H_SCP,
       SPI1_SS3_F2H_SCP,
       TX_CLKPF,
       USER_MSS_GPIO_RESET_N,
       USER_MSS_RESET_N,
       XCLK_FAB,
       CLK_BASE,
       CLK_MDDR_APB,
       F_ARADDR_HADDR1,
       F_ARBURST_HTRANS1,
       F_ARID_HSEL1,
       F_ARLEN_HBURST1,
       F_ARLOCK_HMASTLOCK1,
       F_ARSIZE_HSIZE1,
       F_ARVALID_HWRITE1,
       F_AWADDR_HADDR0,
       F_AWBURST_HTRANS0,
       F_AWID_HSEL0,
       F_AWLEN_HBURST0,
       F_AWLOCK_HMASTLOCK0,
       F_AWSIZE_HSIZE0,
       F_AWVALID_HWRITE0,
       F_BREADY,
       F_RMW_AXI,
       F_RREADY,
       F_WDATA_HWDATA01,
       F_WID_HREADY01,
       F_WLAST,
       F_WSTRB,
       F_WVALID,
       FPGA_MDDR_ARESET_N,
       MDDR_FABRIC_PADDR,
       MDDR_FABRIC_PENABLE,
       MDDR_FABRIC_PSEL,
       MDDR_FABRIC_PWDATA,
       MDDR_FABRIC_PWRITE,
       PRESET_N,
       CAN_RXBUS_USBA_DATA1_MGPIO3A_IN,
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN,
       CAN_TXBUS_USBA_DATA0_MGPIO2A_IN,
       DM_IN,
       DRAM_DQ_IN,
       DRAM_DQS_IN,
       DRAM_FIFO_WE_IN,
       I2C0_SCL_USBC_DATA1_MGPIO31B_IN,
       I2C0_SDA_USBC_DATA0_MGPIO30B_IN,
       I2C1_SCL_USBA_DATA4_MGPIO1A_IN,
       I2C1_SDA_USBA_DATA3_MGPIO0A_IN,
       MMUART0_CTS_USBC_DATA7_MGPIO19B_IN,
       MMUART0_DCD_MGPIO22B_IN,
       MMUART0_DSR_MGPIO20B_IN,
       MMUART0_DTR_USBC_DATA6_MGPIO18B_IN,
       MMUART0_RI_MGPIO21B_IN,
       MMUART0_RTS_USBC_DATA5_MGPIO17B_IN,
       MMUART0_RXD_USBC_STP_MGPIO28B_IN,
       MMUART0_SCK_USBC_NXT_MGPIO29B_IN,
       MMUART0_TXD_USBC_DIR_MGPIO27B_IN,
       MMUART1_RXD_USBC_DATA3_MGPIO26B_IN,
       MMUART1_SCK_USBC_DATA4_MGPIO25B_IN,
       MMUART1_TXD_USBC_DATA2_MGPIO24B_IN,
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN,
       RGMII_MDC_RMII_MDC_IN,
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN,
       RGMII_RX_CLK_IN,
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN,
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN,
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN,
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN,
       RGMII_RXD3_USBB_DATA4_IN,
       RGMII_TX_CLK_IN,
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN,
       RGMII_TXD0_RMII_TXD0_USBB_DIR_IN,
       RGMII_TXD1_RMII_TXD1_USBB_STP_IN,
       RGMII_TXD2_USBB_DATA5_IN,
       RGMII_TXD3_USBB_DATA6_IN,
       SPI0_SCK_USBA_XCLK_IN,
       SPI0_SDI_USBA_DIR_MGPIO5A_IN,
       SPI0_SDO_USBA_STP_MGPIO6A_IN,
       SPI0_SS0_USBA_NXT_MGPIO7A_IN,
       SPI0_SS1_USBA_DATA5_MGPIO8A_IN,
       SPI0_SS2_USBA_DATA6_MGPIO9A_IN,
       SPI0_SS3_USBA_DATA7_MGPIO10A_IN,
       SPI1_SCK_IN,
       SPI1_SDI_MGPIO11A_IN,
       SPI1_SDO_MGPIO12A_IN,
       SPI1_SS0_MGPIO13A_IN,
       SPI1_SS1_MGPIO14A_IN,
       SPI1_SS2_MGPIO15A_IN,
       SPI1_SS3_MGPIO16A_IN,
       SPI1_SS4_MGPIO17A_IN,
       SPI1_SS5_MGPIO18A_IN,
       SPI1_SS6_MGPIO23A_IN,
       SPI1_SS7_MGPIO24A_IN,
       USBC_XCLK_IN,
       CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT,
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT,
       CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT,
       DRAM_ADDR,
       DRAM_BA,
       DRAM_CASN,
       DRAM_CKE,
       DRAM_CLK,
       DRAM_CSN,
       DRAM_DM_RDQS_OUT,
       DRAM_DQ_OUT,
       DRAM_DQS_OUT,
       DRAM_FIFO_WE_OUT,
       DRAM_ODT,
       DRAM_RASN,
       DRAM_RSTN,
       DRAM_WEN,
       I2C0_SCL_USBC_DATA1_MGPIO31B_OUT,
       I2C0_SDA_USBC_DATA0_MGPIO30B_OUT,
       I2C1_SCL_USBA_DATA4_MGPIO1A_OUT,
       I2C1_SDA_USBA_DATA3_MGPIO0A_OUT,
       MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT,
       MMUART0_DCD_MGPIO22B_OUT,
       MMUART0_DSR_MGPIO20B_OUT,
       MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT,
       MMUART0_RI_MGPIO21B_OUT,
       MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT,
       MMUART0_RXD_USBC_STP_MGPIO28B_OUT,
       MMUART0_SCK_USBC_NXT_MGPIO29B_OUT,
       MMUART0_TXD_USBC_DIR_MGPIO27B_OUT,
       MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT,
       MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT,
       MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT,
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT,
       RGMII_MDC_RMII_MDC_OUT,
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT,
       RGMII_RX_CLK_OUT,
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT,
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT,
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT,
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT,
       RGMII_RXD3_USBB_DATA4_OUT,
       RGMII_TX_CLK_OUT,
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT,
       RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT,
       RGMII_TXD1_RMII_TXD1_USBB_STP_OUT,
       RGMII_TXD2_USBB_DATA5_OUT,
       RGMII_TXD3_USBB_DATA6_OUT,
       SPI0_SCK_USBA_XCLK_OUT,
       SPI0_SDI_USBA_DIR_MGPIO5A_OUT,
       SPI0_SDO_USBA_STP_MGPIO6A_OUT,
       SPI0_SS0_USBA_NXT_MGPIO7A_OUT,
       SPI0_SS1_USBA_DATA5_MGPIO8A_OUT,
       SPI0_SS2_USBA_DATA6_MGPIO9A_OUT,
       SPI0_SS3_USBA_DATA7_MGPIO10A_OUT,
       SPI1_SCK_OUT,
       SPI1_SDI_MGPIO11A_OUT,
       SPI1_SDO_MGPIO12A_OUT,
       SPI1_SS0_MGPIO13A_OUT,
       SPI1_SS1_MGPIO14A_OUT,
       SPI1_SS2_MGPIO15A_OUT,
       SPI1_SS3_MGPIO16A_OUT,
       SPI1_SS4_MGPIO17A_OUT,
       SPI1_SS5_MGPIO18A_OUT,
       SPI1_SS6_MGPIO23A_OUT,
       SPI1_SS7_MGPIO24A_OUT,
       USBC_XCLK_OUT,
       CAN_RXBUS_USBA_DATA1_MGPIO3A_OE,
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE,
       CAN_TXBUS_USBA_DATA0_MGPIO2A_OE,
       DM_OE,
       DRAM_DQ_OE,
       DRAM_DQS_OE,
       I2C0_SCL_USBC_DATA1_MGPIO31B_OE,
       I2C0_SDA_USBC_DATA0_MGPIO30B_OE,
       I2C1_SCL_USBA_DATA4_MGPIO1A_OE,
       I2C1_SDA_USBA_DATA3_MGPIO0A_OE,
       MMUART0_CTS_USBC_DATA7_MGPIO19B_OE,
       MMUART0_DCD_MGPIO22B_OE,
       MMUART0_DSR_MGPIO20B_OE,
       MMUART0_DTR_USBC_DATA6_MGPIO18B_OE,
       MMUART0_RI_MGPIO21B_OE,
       MMUART0_RTS_USBC_DATA5_MGPIO17B_OE,
       MMUART0_RXD_USBC_STP_MGPIO28B_OE,
       MMUART0_SCK_USBC_NXT_MGPIO29B_OE,
       MMUART0_TXD_USBC_DIR_MGPIO27B_OE,
       MMUART1_RXD_USBC_DATA3_MGPIO26B_OE,
       MMUART1_SCK_USBC_DATA4_MGPIO25B_OE,
       MMUART1_TXD_USBC_DATA2_MGPIO24B_OE,
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE,
       RGMII_MDC_RMII_MDC_OE,
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE,
       RGMII_RX_CLK_OE,
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE,
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE,
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE,
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE,
       RGMII_RXD3_USBB_DATA4_OE,
       RGMII_TX_CLK_OE,
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE,
       RGMII_TXD0_RMII_TXD0_USBB_DIR_OE,
       RGMII_TXD1_RMII_TXD1_USBB_STP_OE,
       RGMII_TXD2_USBB_DATA5_OE,
       RGMII_TXD3_USBB_DATA6_OE,
       SPI0_SCK_USBA_XCLK_OE,
       SPI0_SDI_USBA_DIR_MGPIO5A_OE,
       SPI0_SDO_USBA_STP_MGPIO6A_OE,
       SPI0_SS0_USBA_NXT_MGPIO7A_OE,
       SPI0_SS1_USBA_DATA5_MGPIO8A_OE,
       SPI0_SS2_USBA_DATA6_MGPIO9A_OE,
       SPI0_SS3_USBA_DATA7_MGPIO10A_OE,
       SPI1_SCK_OE,
       SPI1_SDI_MGPIO11A_OE,
       SPI1_SDO_MGPIO12A_OE,
       SPI1_SS0_MGPIO13A_OE,
       SPI1_SS1_MGPIO14A_OE,
       SPI1_SS2_MGPIO15A_OE,
       SPI1_SS3_MGPIO16A_OE,
       SPI1_SS4_MGPIO17A_OE,
       SPI1_SS5_MGPIO18A_OE,
       SPI1_SS6_MGPIO23A_OE,
       SPI1_SS7_MGPIO24A_OE,
       USBC_XCLK_OE
    );
output CAN_RXBUS_MGPIO3A_H2F_A;
output CAN_RXBUS_MGPIO3A_H2F_B;
output CAN_TX_EBL_MGPIO4A_H2F_A;
output CAN_TX_EBL_MGPIO4A_H2F_B;
output CAN_TXBUS_MGPIO2A_H2F_A;
output CAN_TXBUS_MGPIO2A_H2F_B;
output CLK_CONFIG_APB;
output COMMS_INT;
output CONFIG_PRESET_N;
output [7:0] EDAC_ERROR;
output [31:0] F_FM0_RDATA;
output F_FM0_READYOUT;
output F_FM0_RESP;
output [31:0] F_HM0_ADDR;
output F_HM0_ENABLE;
output F_HM0_SEL;
output [1:0] F_HM0_SIZE;
output F_HM0_TRANS1;
output [31:0] F_HM0_WDATA;
output F_HM0_WRITE;
output FAB_CHRGVBUS;
output FAB_DISCHRGVBUS;
output FAB_DMPULLDOWN;
output FAB_DPPULLDOWN;
output FAB_DRVVBUS;
output FAB_IDPULLUP;
output [1:0] FAB_OPMODE;
output FAB_SUSPENDM;
output FAB_TERMSEL;
output FAB_TXVALID;
output [3:0] FAB_VCONTROL;
output FAB_VCONTROLLOADM;
output [1:0] FAB_XCVRSEL;
output [7:0] FAB_XDATAOUT;
output FACC_GLMUX_SEL;
output [1:0] FIC32_0_MASTER;
output [1:0] FIC32_1_MASTER;
output FPGA_RESET_N;
output GTX_CLK;
output [15:0] H2F_INTERRUPT;
output H2F_NMI;
output H2FCALIB;
output I2C0_SCL_MGPIO31B_H2F_A;
output I2C0_SCL_MGPIO31B_H2F_B;
output I2C0_SDA_MGPIO30B_H2F_A;
output I2C0_SDA_MGPIO30B_H2F_B;
output I2C1_SCL_MGPIO1A_H2F_A;
output I2C1_SCL_MGPIO1A_H2F_B;
output I2C1_SDA_MGPIO0A_H2F_A;
output I2C1_SDA_MGPIO0A_H2F_B;
output MDCF;
output MDOENF;
output MDOF;
output MMUART0_CTS_MGPIO19B_H2F_A;
output MMUART0_CTS_MGPIO19B_H2F_B;
output MMUART0_DCD_MGPIO22B_H2F_A;
output MMUART0_DCD_MGPIO22B_H2F_B;
output MMUART0_DSR_MGPIO20B_H2F_A;
output MMUART0_DSR_MGPIO20B_H2F_B;
output MMUART0_DTR_MGPIO18B_H2F_A;
output MMUART0_DTR_MGPIO18B_H2F_B;
output MMUART0_RI_MGPIO21B_H2F_A;
output MMUART0_RI_MGPIO21B_H2F_B;
output MMUART0_RTS_MGPIO17B_H2F_A;
output MMUART0_RTS_MGPIO17B_H2F_B;
output MMUART0_RXD_MGPIO28B_H2F_A;
output MMUART0_RXD_MGPIO28B_H2F_B;
output MMUART0_SCK_MGPIO29B_H2F_A;
output MMUART0_SCK_MGPIO29B_H2F_B;
output MMUART0_TXD_MGPIO27B_H2F_A;
output MMUART0_TXD_MGPIO27B_H2F_B;
output MMUART1_DTR_MGPIO12B_H2F_A;
output MMUART1_RTS_MGPIO11B_H2F_A;
output MMUART1_RTS_MGPIO11B_H2F_B;
output MMUART1_RXD_MGPIO26B_H2F_A;
output MMUART1_RXD_MGPIO26B_H2F_B;
output MMUART1_SCK_MGPIO25B_H2F_A;
output MMUART1_SCK_MGPIO25B_H2F_B;
output MMUART1_TXD_MGPIO24B_H2F_A;
output MMUART1_TXD_MGPIO24B_H2F_B;
output MPLL_LOCK;
output [15:2] PER2_FABRIC_PADDR;
output PER2_FABRIC_PENABLE;
output PER2_FABRIC_PSEL;
output [31:0] PER2_FABRIC_PWDATA;
output PER2_FABRIC_PWRITE;
output RTC_MATCH;
output SLEEPDEEP;
output SLEEPHOLDACK;
output SLEEPING;
output SMBALERT_NO0;
output SMBALERT_NO1;
output SMBSUS_NO0;
output SMBSUS_NO1;
output SPI0_CLK_OUT;
output SPI0_SDI_MGPIO5A_H2F_A;
output SPI0_SDI_MGPIO5A_H2F_B;
output SPI0_SDO_MGPIO6A_H2F_A;
output SPI0_SDO_MGPIO6A_H2F_B;
output SPI0_SS0_MGPIO7A_H2F_A;
output SPI0_SS0_MGPIO7A_H2F_B;
output SPI0_SS1_MGPIO8A_H2F_A;
output SPI0_SS1_MGPIO8A_H2F_B;
output SPI0_SS2_MGPIO9A_H2F_A;
output SPI0_SS2_MGPIO9A_H2F_B;
output SPI0_SS3_MGPIO10A_H2F_A;
output SPI0_SS3_MGPIO10A_H2F_B;
output SPI0_SS4_MGPIO19A_H2F_A;
output SPI0_SS5_MGPIO20A_H2F_A;
output SPI0_SS6_MGPIO21A_H2F_A;
output SPI0_SS7_MGPIO22A_H2F_A;
output SPI1_CLK_OUT;
output SPI1_SDI_MGPIO11A_H2F_A;
output SPI1_SDI_MGPIO11A_H2F_B;
output SPI1_SDO_MGPIO12A_H2F_A;
output SPI1_SDO_MGPIO12A_H2F_B;
output SPI1_SS0_MGPIO13A_H2F_A;
output SPI1_SS0_MGPIO13A_H2F_B;
output SPI1_SS1_MGPIO14A_H2F_A;
output SPI1_SS1_MGPIO14A_H2F_B;
output SPI1_SS2_MGPIO15A_H2F_A;
output SPI1_SS2_MGPIO15A_H2F_B;
output SPI1_SS3_MGPIO16A_H2F_A;
output SPI1_SS3_MGPIO16A_H2F_B;
output SPI1_SS4_MGPIO17A_H2F_A;
output SPI1_SS5_MGPIO18A_H2F_A;
output SPI1_SS6_MGPIO23A_H2F_A;
output SPI1_SS7_MGPIO24A_H2F_A;
output [9:0] TCGF;
output TRACECLK;
output [3:0] TRACEDATA;
output TX_CLK;
output TX_ENF;
output TX_ERRF;
output TXCTL_EN_RIF;
output [3:0] TXD_RIF;
output [7:0] TXDF;
output TXEV;
output WDOGTIMEOUT;
output F_ARREADY_HREADYOUT1;
output F_AWREADY_HREADYOUT0;
output [3:0] F_BID;
output [1:0] F_BRESP_HRESP0;
output F_BVALID;
output [63:0] F_RDATA_HRDATA01;
output [3:0] F_RID;
output F_RLAST;
output [1:0] F_RRESP_HRESP1;
output F_RVALID;
output F_WREADY;
output [15:0] MDDR_FABRIC_PRDATA;
output MDDR_FABRIC_PREADY;
output MDDR_FABRIC_PSLVERR;
input  CAN_RXBUS_F2H_SCP;
input  CAN_TX_EBL_F2H_SCP;
input  CAN_TXBUS_F2H_SCP;
input  COLF;
input  CRSF;
input  [1:0] F2_DMAREADY;
input  [15:0] F2H_INTERRUPT;
input  F2HCALIB;
input  [1:0] F_DMAREADY;
input  [31:0] F_FM0_ADDR;
input  F_FM0_ENABLE;
input  F_FM0_MASTLOCK;
input  F_FM0_READY;
input  F_FM0_SEL;
input  [1:0] F_FM0_SIZE;
input  F_FM0_TRANS1;
input  [31:0] F_FM0_WDATA;
input  F_FM0_WRITE;
input  [31:0] F_HM0_RDATA;
input  F_HM0_READY;
input  F_HM0_RESP;
input  FAB_AVALID;
input  FAB_HOSTDISCON;
input  FAB_IDDIG;
input  [1:0] FAB_LINESTATE;
input  FAB_M3_RESET_N;
input  FAB_PLL_LOCK;
input  FAB_RXACTIVE;
input  FAB_RXERROR;
input  FAB_RXVALID;
input  FAB_RXVALIDH;
input  FAB_SESSEND;
input  FAB_TXREADY;
input  FAB_VBUSVALID;
input  [7:0] FAB_VSTATUS;
input  [7:0] FAB_XDATAIN;
input  GTX_CLKPF;
input  I2C0_BCLK;
input  I2C0_SCL_F2H_SCP;
input  I2C0_SDA_F2H_SCP;
input  I2C1_BCLK;
input  I2C1_SCL_F2H_SCP;
input  I2C1_SDA_F2H_SCP;
input  MDIF;
input  MGPIO0A_F2H_GPIN;
input  MGPIO10A_F2H_GPIN;
input  MGPIO11A_F2H_GPIN;
input  MGPIO11B_F2H_GPIN;
input  MGPIO12A_F2H_GPIN;
input  MGPIO13A_F2H_GPIN;
input  MGPIO14A_F2H_GPIN;
input  MGPIO15A_F2H_GPIN;
input  MGPIO16A_F2H_GPIN;
input  MGPIO17B_F2H_GPIN;
input  MGPIO18B_F2H_GPIN;
input  MGPIO19B_F2H_GPIN;
input  MGPIO1A_F2H_GPIN;
input  MGPIO20B_F2H_GPIN;
input  MGPIO21B_F2H_GPIN;
input  MGPIO22B_F2H_GPIN;
input  MGPIO24B_F2H_GPIN;
input  MGPIO25B_F2H_GPIN;
input  MGPIO26B_F2H_GPIN;
input  MGPIO27B_F2H_GPIN;
input  MGPIO28B_F2H_GPIN;
input  MGPIO29B_F2H_GPIN;
input  MGPIO2A_F2H_GPIN;
input  MGPIO30B_F2H_GPIN;
input  MGPIO31B_F2H_GPIN;
input  MGPIO3A_F2H_GPIN;
input  MGPIO4A_F2H_GPIN;
input  MGPIO5A_F2H_GPIN;
input  MGPIO6A_F2H_GPIN;
input  MGPIO7A_F2H_GPIN;
input  MGPIO8A_F2H_GPIN;
input  MGPIO9A_F2H_GPIN;
input  MMUART0_CTS_F2H_SCP;
input  MMUART0_DCD_F2H_SCP;
input  MMUART0_DSR_F2H_SCP;
input  MMUART0_DTR_F2H_SCP;
input  MMUART0_RI_F2H_SCP;
input  MMUART0_RTS_F2H_SCP;
input  MMUART0_RXD_F2H_SCP;
input  MMUART0_SCK_F2H_SCP;
input  MMUART0_TXD_F2H_SCP;
input  MMUART1_CTS_F2H_SCP;
input  MMUART1_DCD_F2H_SCP;
input  MMUART1_DSR_F2H_SCP;
input  MMUART1_RI_F2H_SCP;
input  MMUART1_RTS_F2H_SCP;
input  MMUART1_RXD_F2H_SCP;
input  MMUART1_SCK_F2H_SCP;
input  MMUART1_TXD_F2H_SCP;
input  [31:0] PER2_FABRIC_PRDATA;
input  PER2_FABRIC_PREADY;
input  PER2_FABRIC_PSLVERR;
input  [9:0] RCGF;
input  RX_CLKPF;
input  RX_DVF;
input  RX_ERRF;
input  RX_EV;
input  [7:0] RXDF;
input  SLEEPHOLDREQ;
input  SMBALERT_NI0;
input  SMBALERT_NI1;
input  SMBSUS_NI0;
input  SMBSUS_NI1;
input  SPI0_CLK_IN;
input  SPI0_SDI_F2H_SCP;
input  SPI0_SDO_F2H_SCP;
input  SPI0_SS0_F2H_SCP;
input  SPI0_SS1_F2H_SCP;
input  SPI0_SS2_F2H_SCP;
input  SPI0_SS3_F2H_SCP;
input  SPI1_CLK_IN;
input  SPI1_SDI_F2H_SCP;
input  SPI1_SDO_F2H_SCP;
input  SPI1_SS0_F2H_SCP;
input  SPI1_SS1_F2H_SCP;
input  SPI1_SS2_F2H_SCP;
input  SPI1_SS3_F2H_SCP;
input  TX_CLKPF;
input  USER_MSS_GPIO_RESET_N;
input  USER_MSS_RESET_N;
input  XCLK_FAB;
input  CLK_BASE;
input  CLK_MDDR_APB;
input  [31:0] F_ARADDR_HADDR1;
input  [1:0] F_ARBURST_HTRANS1;
input  [3:0] F_ARID_HSEL1;
input  [3:0] F_ARLEN_HBURST1;
input  [1:0] F_ARLOCK_HMASTLOCK1;
input  [1:0] F_ARSIZE_HSIZE1;
input  F_ARVALID_HWRITE1;
input  [31:0] F_AWADDR_HADDR0;
input  [1:0] F_AWBURST_HTRANS0;
input  [3:0] F_AWID_HSEL0;
input  [3:0] F_AWLEN_HBURST0;
input  [1:0] F_AWLOCK_HMASTLOCK0;
input  [1:0] F_AWSIZE_HSIZE0;
input  F_AWVALID_HWRITE0;
input  F_BREADY;
input  F_RMW_AXI;
input  F_RREADY;
input  [63:0] F_WDATA_HWDATA01;
input  [3:0] F_WID_HREADY01;
input  F_WLAST;
input  [7:0] F_WSTRB;
input  F_WVALID;
input  FPGA_MDDR_ARESET_N;
input  [10:2] MDDR_FABRIC_PADDR;
input  MDDR_FABRIC_PENABLE;
input  MDDR_FABRIC_PSEL;
input  [15:0] MDDR_FABRIC_PWDATA;
input  MDDR_FABRIC_PWRITE;
input  PRESET_N;
input  CAN_RXBUS_USBA_DATA1_MGPIO3A_IN;
input  CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN;
input  CAN_TXBUS_USBA_DATA0_MGPIO2A_IN;
input  [2:0] DM_IN;
input  [17:0] DRAM_DQ_IN;
input  [2:0] DRAM_DQS_IN;
input  [1:0] DRAM_FIFO_WE_IN;
input  I2C0_SCL_USBC_DATA1_MGPIO31B_IN;
input  I2C0_SDA_USBC_DATA0_MGPIO30B_IN;
input  I2C1_SCL_USBA_DATA4_MGPIO1A_IN;
input  I2C1_SDA_USBA_DATA3_MGPIO0A_IN;
input  MMUART0_CTS_USBC_DATA7_MGPIO19B_IN;
input  MMUART0_DCD_MGPIO22B_IN;
input  MMUART0_DSR_MGPIO20B_IN;
input  MMUART0_DTR_USBC_DATA6_MGPIO18B_IN;
input  MMUART0_RI_MGPIO21B_IN;
input  MMUART0_RTS_USBC_DATA5_MGPIO17B_IN;
input  MMUART0_RXD_USBC_STP_MGPIO28B_IN;
input  MMUART0_SCK_USBC_NXT_MGPIO29B_IN;
input  MMUART0_TXD_USBC_DIR_MGPIO27B_IN;
input  MMUART1_RXD_USBC_DATA3_MGPIO26B_IN;
input  MMUART1_SCK_USBC_DATA4_MGPIO25B_IN;
input  MMUART1_TXD_USBC_DATA2_MGPIO24B_IN;
input  RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN;
input  RGMII_MDC_RMII_MDC_IN;
input  RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN;
input  RGMII_RX_CLK_IN;
input  RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN;
input  RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN;
input  RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN;
input  RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN;
input  RGMII_RXD3_USBB_DATA4_IN;
input  RGMII_TX_CLK_IN;
input  RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN;
input  RGMII_TXD0_RMII_TXD0_USBB_DIR_IN;
input  RGMII_TXD1_RMII_TXD1_USBB_STP_IN;
input  RGMII_TXD2_USBB_DATA5_IN;
input  RGMII_TXD3_USBB_DATA6_IN;
input  SPI0_SCK_USBA_XCLK_IN;
input  SPI0_SDI_USBA_DIR_MGPIO5A_IN;
input  SPI0_SDO_USBA_STP_MGPIO6A_IN;
input  SPI0_SS0_USBA_NXT_MGPIO7A_IN;
input  SPI0_SS1_USBA_DATA5_MGPIO8A_IN;
input  SPI0_SS2_USBA_DATA6_MGPIO9A_IN;
input  SPI0_SS3_USBA_DATA7_MGPIO10A_IN;
input  SPI1_SCK_IN;
input  SPI1_SDI_MGPIO11A_IN;
input  SPI1_SDO_MGPIO12A_IN;
input  SPI1_SS0_MGPIO13A_IN;
input  SPI1_SS1_MGPIO14A_IN;
input  SPI1_SS2_MGPIO15A_IN;
input  SPI1_SS3_MGPIO16A_IN;
input  SPI1_SS4_MGPIO17A_IN;
input  SPI1_SS5_MGPIO18A_IN;
input  SPI1_SS6_MGPIO23A_IN;
input  SPI1_SS7_MGPIO24A_IN;
input  USBC_XCLK_IN;
output CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT;
output CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT;
output CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT;
output [15:0] DRAM_ADDR;
output [2:0] DRAM_BA;
output DRAM_CASN;
output DRAM_CKE;
output DRAM_CLK;
output DRAM_CSN;
output [2:0] DRAM_DM_RDQS_OUT;
output [17:0] DRAM_DQ_OUT;
output [2:0] DRAM_DQS_OUT;
output [1:0] DRAM_FIFO_WE_OUT;
output DRAM_ODT;
output DRAM_RASN;
output DRAM_RSTN;
output DRAM_WEN;
output I2C0_SCL_USBC_DATA1_MGPIO31B_OUT;
output I2C0_SDA_USBC_DATA0_MGPIO30B_OUT;
output I2C1_SCL_USBA_DATA4_MGPIO1A_OUT;
output I2C1_SDA_USBA_DATA3_MGPIO0A_OUT;
output MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT;
output MMUART0_DCD_MGPIO22B_OUT;
output MMUART0_DSR_MGPIO20B_OUT;
output MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT;
output MMUART0_RI_MGPIO21B_OUT;
output MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT;
output MMUART0_RXD_USBC_STP_MGPIO28B_OUT;
output MMUART0_SCK_USBC_NXT_MGPIO29B_OUT;
output MMUART0_TXD_USBC_DIR_MGPIO27B_OUT;
output MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT;
output MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT;
output MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT;
output RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT;
output RGMII_MDC_RMII_MDC_OUT;
output RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT;
output RGMII_RX_CLK_OUT;
output RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT;
output RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT;
output RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT;
output RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT;
output RGMII_RXD3_USBB_DATA4_OUT;
output RGMII_TX_CLK_OUT;
output RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT;
output RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT;
output RGMII_TXD1_RMII_TXD1_USBB_STP_OUT;
output RGMII_TXD2_USBB_DATA5_OUT;
output RGMII_TXD3_USBB_DATA6_OUT;
output SPI0_SCK_USBA_XCLK_OUT;
output SPI0_SDI_USBA_DIR_MGPIO5A_OUT;
output SPI0_SDO_USBA_STP_MGPIO6A_OUT;
output SPI0_SS0_USBA_NXT_MGPIO7A_OUT;
output SPI0_SS1_USBA_DATA5_MGPIO8A_OUT;
output SPI0_SS2_USBA_DATA6_MGPIO9A_OUT;
output SPI0_SS3_USBA_DATA7_MGPIO10A_OUT;
output SPI1_SCK_OUT;
output SPI1_SDI_MGPIO11A_OUT;
output SPI1_SDO_MGPIO12A_OUT;
output SPI1_SS0_MGPIO13A_OUT;
output SPI1_SS1_MGPIO14A_OUT;
output SPI1_SS2_MGPIO15A_OUT;
output SPI1_SS3_MGPIO16A_OUT;
output SPI1_SS4_MGPIO17A_OUT;
output SPI1_SS5_MGPIO18A_OUT;
output SPI1_SS6_MGPIO23A_OUT;
output SPI1_SS7_MGPIO24A_OUT;
output USBC_XCLK_OUT;
output CAN_RXBUS_USBA_DATA1_MGPIO3A_OE;
output CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE;
output CAN_TXBUS_USBA_DATA0_MGPIO2A_OE;
output [2:0] DM_OE;
output [17:0] DRAM_DQ_OE;
output [2:0] DRAM_DQS_OE;
output I2C0_SCL_USBC_DATA1_MGPIO31B_OE;
output I2C0_SDA_USBC_DATA0_MGPIO30B_OE;
output I2C1_SCL_USBA_DATA4_MGPIO1A_OE;
output I2C1_SDA_USBA_DATA3_MGPIO0A_OE;
output MMUART0_CTS_USBC_DATA7_MGPIO19B_OE;
output MMUART0_DCD_MGPIO22B_OE;
output MMUART0_DSR_MGPIO20B_OE;
output MMUART0_DTR_USBC_DATA6_MGPIO18B_OE;
output MMUART0_RI_MGPIO21B_OE;
output MMUART0_RTS_USBC_DATA5_MGPIO17B_OE;
output MMUART0_RXD_USBC_STP_MGPIO28B_OE;
output MMUART0_SCK_USBC_NXT_MGPIO29B_OE;
output MMUART0_TXD_USBC_DIR_MGPIO27B_OE;
output MMUART1_RXD_USBC_DATA3_MGPIO26B_OE;
output MMUART1_SCK_USBC_DATA4_MGPIO25B_OE;
output MMUART1_TXD_USBC_DATA2_MGPIO24B_OE;
output RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE;
output RGMII_MDC_RMII_MDC_OE;
output RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE;
output RGMII_RX_CLK_OE;
output RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE;
output RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE;
output RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE;
output RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE;
output RGMII_RXD3_USBB_DATA4_OE;
output RGMII_TX_CLK_OE;
output RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE;
output RGMII_TXD0_RMII_TXD0_USBB_DIR_OE;
output RGMII_TXD1_RMII_TXD1_USBB_STP_OE;
output RGMII_TXD2_USBB_DATA5_OE;
output RGMII_TXD3_USBB_DATA6_OE;
output SPI0_SCK_USBA_XCLK_OE;
output SPI0_SDI_USBA_DIR_MGPIO5A_OE;
output SPI0_SDO_USBA_STP_MGPIO6A_OE;
output SPI0_SS0_USBA_NXT_MGPIO7A_OE;
output SPI0_SS1_USBA_DATA5_MGPIO8A_OE;
output SPI0_SS2_USBA_DATA6_MGPIO9A_OE;
output SPI0_SS3_USBA_DATA7_MGPIO10A_OE;
output SPI1_SCK_OE;
output SPI1_SDI_MGPIO11A_OE;
output SPI1_SDO_MGPIO12A_OE;
output SPI1_SS0_MGPIO13A_OE;
output SPI1_SS1_MGPIO14A_OE;
output SPI1_SS2_MGPIO15A_OE;
output SPI1_SS3_MGPIO16A_OE;
output SPI1_SS4_MGPIO17A_OE;
output SPI1_SS5_MGPIO18A_OE;
output SPI1_SS6_MGPIO23A_OE;
output SPI1_SS7_MGPIO24A_OE;
output USBC_XCLK_OE;

    parameter INIT = 'h0 ;
    parameter ACT_UBITS = 'hFFFFFFFFFFFFFF ;
    parameter MEMORYFILE = "" ;
    parameter RTC_MAIN_XTL_FREQ = 0.0 ;
    parameter RTC_MAIN_XTL_MODE = "1" ;
    parameter DDR_CLK_FREQ = 0.0 ;
    
endmodule


module SF2Project_MSS(
       MDDR_DQS,
       MDDR_DQS_N,
       MAC_MII_RXD,
       MAC_MII_TXD,
       MDDR_ADDR,
       MDDR_BA,
       MDDR_DM_RDQS,
       MDDR_DQ,
       USB_ULPI_DATA,
       MDDR_CLK,
       MDDR_CLK_N,
       MCCC_CLK_BASE,
       MAC_MII_TX_CLK,
       MAC_MII_RX_ER,
       MAC_MII_RX_DV,
       MAC_MII_RX_CLK,
       MAC_MII_CRS,
       MAC_MII_COL,
       MAC_MII_TX_ER,
       MAC_MII_TX_EN,
       I2C_0_SCL,
       I2C_0_SDA,
       I2C_1_SCL,
       I2C_1_SDA,
       MDDR_CAS_N,
       MDDR_CKE,
       MDDR_CS_N,
       MDDR_DQS_TMATCH_0_IN,
       MDDR_DQS_TMATCH_0_OUT,
       MDDR_ODT,
       MDDR_RAS_N,
       MDDR_RESET_N,
       MDDR_WE_N,
       MMUART_0_RXD,
       MMUART_0_TXD,
       MMUART_1_RXD,
       MMUART_1_TXD,
       SPI_0_CLK,
       SPI_0_DI,
       SPI_0_DO,
       SPI_0_SS0,
       SPI_1_CLK,
       SPI_1_DI,
       SPI_1_DO,
       SPI_1_SS0,
       USB_ULPI_DIR,
       USB_ULPI_NXT,
       USB_ULPI_STP,
       USB_ULPI_XCLK
    );
inout  [1:0] MDDR_DQS;
inout  [1:0] MDDR_DQS_N;
input  [3:0] MAC_MII_RXD;
output [3:0] MAC_MII_TXD;
output [15:0] MDDR_ADDR;
output [2:0] MDDR_BA;
inout  [1:0] MDDR_DM_RDQS;
inout  [15:0] MDDR_DQ;
inout  [7:0] USB_ULPI_DATA;
output MDDR_CLK;
output MDDR_CLK_N;
input  MCCC_CLK_BASE;
input  MAC_MII_TX_CLK;
input  MAC_MII_RX_ER;
input  MAC_MII_RX_DV;
input  MAC_MII_RX_CLK;
input  MAC_MII_CRS;
input  MAC_MII_COL;
output MAC_MII_TX_ER;
output MAC_MII_TX_EN;
inout  I2C_0_SCL;
inout  I2C_0_SDA;
inout  I2C_1_SCL;
inout  I2C_1_SDA;
output MDDR_CAS_N;
output MDDR_CKE;
output MDDR_CS_N;
input  MDDR_DQS_TMATCH_0_IN;
output MDDR_DQS_TMATCH_0_OUT;
output MDDR_ODT;
output MDDR_RAS_N;
output MDDR_RESET_N;
output MDDR_WE_N;
input  MMUART_0_RXD;
output MMUART_0_TXD;
input  MMUART_1_RXD;
output MMUART_1_TXD;
inout  SPI_0_CLK;
input  SPI_0_DI;
output SPI_0_DO;
inout  SPI_0_SS0;
inout  SPI_1_CLK;
input  SPI_1_DI;
output SPI_1_DO;
inout  SPI_1_SS0;
input  USB_ULPI_DIR;
input  USB_ULPI_NXT;
output USB_ULPI_STP;
input  USB_ULPI_XCLK;

    wire [1:0] DRAM_FIFO_WE_OUT_net_0;
    wire [17:0] DRAM_DQ_OUT_net_0;
    wire [17:0] DRAM_DQ_OE_net_0;
    wire [2:0] DRAM_DM_RDQS_OUT_net_0;
    wire [2:0] DM_OE_net_0;
    wire [2:0] DRAM_BA_net_0;
    wire [15:0] DRAM_ADDR_net_0;
    wire [7:0] EDAC_ERROR;
    wire [31:0] F_FM0_RDATA;
    wire [31:0] F_HM0_ADDR;
    wire [1:0] F_HM0_SIZE;
    wire [31:0] F_HM0_WDATA;
    wire [1:0] FAB_OPMODE;
    wire [3:0] FAB_VCONTROL;
    wire [1:0] FAB_XCVRSEL;
    wire [7:0] FAB_XDATAOUT;
    wire [1:0] FIC32_0_MASTER;
    wire [1:0] FIC32_1_MASTER;
    wire [15:0] H2F_INTERRUPT;
    wire [15:2] PER2_FABRIC_PADDR;
    wire [31:0] PER2_FABRIC_PWDATA;
    wire [9:0] TCGF;
    wire [3:0] TRACEDATA;
    wire [3:0] TXD_RIF;
    wire [7:4] TXDF_net_0;
    wire [3:0] F_BID;
    wire [1:0] F_BRESP_HRESP0;
    wire [63:0] F_RDATA_HRDATA01;
    wire [3:0] F_RID;
    wire [1:0] F_RRESP_HRESP1;
    wire [15:0] MDDR_FABRIC_PRDATA;
    wire [2:0] DRAM_DQS_OUT_net_0;
    wire [2:0] DRAM_DQS_OE_net_0;
    wire USB_ULPI_XCLK_PAD_Y, 
        MSS_ADLIB_INST_RGMII_TXD1_RMII_TXD1_USBB_STP_OUT, 
        MSS_ADLIB_INST_RGMII_TXD1_RMII_TXD1_USBB_STP_OE, 
        USB_ULPI_NXT_PAD_Y, USB_ULPI_DIR_PAD_Y, USB_ULPI_DATA_7_PAD_Y, 
        MSS_ADLIB_INST_RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT, 
        MSS_ADLIB_INST_RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE, 
        USB_ULPI_DATA_6_PAD_Y, 
        MSS_ADLIB_INST_RGMII_TXD3_USBB_DATA6_OUT, 
        MSS_ADLIB_INST_RGMII_TXD3_USBB_DATA6_OE, USB_ULPI_DATA_5_PAD_Y, 
        MSS_ADLIB_INST_RGMII_TXD2_USBB_DATA5_OUT, 
        MSS_ADLIB_INST_RGMII_TXD2_USBB_DATA5_OE, USB_ULPI_DATA_4_PAD_Y, 
        MSS_ADLIB_INST_RGMII_RXD3_USBB_DATA4_OUT, 
        MSS_ADLIB_INST_RGMII_RXD3_USBB_DATA4_OE, USB_ULPI_DATA_3_PAD_Y, 
        MSS_ADLIB_INST_RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT, 
        MSS_ADLIB_INST_RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE, 
        USB_ULPI_DATA_2_PAD_Y, 
        MSS_ADLIB_INST_RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT, 
        MSS_ADLIB_INST_RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE, 
        USB_ULPI_DATA_1_PAD_Y, 
        MSS_ADLIB_INST_RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT, 
        MSS_ADLIB_INST_RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE, 
        USB_ULPI_DATA_0_PAD_Y, 
        MSS_ADLIB_INST_RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT, 
        MSS_ADLIB_INST_RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE, 
        SPI_1_SS0_PAD_Y, MSS_ADLIB_INST_SPI1_SS0_MGPIO13A_OUT, 
        MSS_ADLIB_INST_SPI1_SS0_MGPIO13A_OE, 
        MSS_ADLIB_INST_SPI1_SDO_MGPIO12A_OUT, 
        MSS_ADLIB_INST_SPI1_SDO_MGPIO12A_OE, SPI_1_DI_PAD_Y, 
        SPI_1_CLK_PAD_Y, MSS_ADLIB_INST_SPI1_SCK_OUT, 
        MSS_ADLIB_INST_SPI1_SCK_OE, SPI_0_SS0_PAD_Y, 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OUT, 
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OE, 
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OUT, 
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OE, SPI_0_DI_PAD_Y, 
        SPI_0_CLK_PAD_Y, MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OUT, 
        MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OE, 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT, 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OE, 
        MMUART_1_RXD_PAD_Y, 
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OUT, 
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OE, 
        MMUART_0_RXD_PAD_Y, MSS_ADLIB_INST_DRAM_WEN, 
        MSS_ADLIB_INST_DRAM_RSTN, MSS_ADLIB_INST_DRAM_RASN, 
        MSS_ADLIB_INST_DRAM_ODT, MDDR_DQS_TMATCH_0_IN_PAD_Y, 
        MDDR_DQ_15_PAD_Y, MDDR_DQ_14_PAD_Y, MDDR_DQ_13_PAD_Y, 
        MDDR_DQ_12_PAD_Y, MDDR_DQ_11_PAD_Y, MDDR_DQ_10_PAD_Y, 
        MDDR_DQ_9_PAD_Y, MDDR_DQ_8_PAD_Y, MDDR_DQ_7_PAD_Y, 
        MDDR_DQ_6_PAD_Y, MDDR_DQ_5_PAD_Y, MDDR_DQ_4_PAD_Y, 
        MDDR_DQ_3_PAD_Y, MDDR_DQ_2_PAD_Y, MDDR_DQ_1_PAD_Y, 
        MDDR_DQ_0_PAD_Y, MDDR_DM_RDQS_1_PAD_Y, MDDR_DM_RDQS_0_PAD_Y, 
        MSS_ADLIB_INST_DRAM_CSN, MSS_ADLIB_INST_DRAM_CKE, 
        MSS_ADLIB_INST_DRAM_CASN, I2C_1_SDA_PAD_Y, 
        MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OUT, 
        MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OE, I2C_1_SCL_PAD_Y, 
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OUT, 
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OE, I2C_0_SDA_PAD_Y, 
        MSS_ADLIB_INST_I2C0_SDA_USBC_DATA0_MGPIO30B_OUT, 
        MSS_ADLIB_INST_I2C0_SDA_USBC_DATA0_MGPIO30B_OE, 
        I2C_0_SCL_PAD_Y, 
        MSS_ADLIB_INST_I2C0_SCL_USBC_DATA1_MGPIO31B_OUT, 
        MSS_ADLIB_INST_I2C0_SCL_USBC_DATA1_MGPIO31B_OE, 
        CAN_RXBUS_MGPIO3A_H2F_A, CAN_RXBUS_MGPIO3A_H2F_B, 
        CAN_TX_EBL_MGPIO4A_H2F_A, CAN_TX_EBL_MGPIO4A_H2F_B, 
        CAN_TXBUS_MGPIO2A_H2F_A, CAN_TXBUS_MGPIO2A_H2F_B, 
        CLK_CONFIG_APB, COMMS_INT, CONFIG_PRESET_N, F_FM0_READYOUT, 
        F_FM0_RESP, F_HM0_ENABLE, F_HM0_SEL, F_HM0_TRANS1, F_HM0_WRITE, 
        FAB_CHRGVBUS, FAB_DISCHRGVBUS, FAB_DMPULLDOWN, FAB_DPPULLDOWN, 
        FAB_DRVVBUS, FAB_IDPULLUP, FAB_SUSPENDM, FAB_TERMSEL, 
        FAB_TXVALID, FAB_VCONTROLLOADM, FACC_GLMUX_SEL, FPGA_RESET_N, 
        GTX_CLK, H2F_NMI, H2FCALIB, I2C0_SCL_MGPIO31B_H2F_A, 
        I2C0_SCL_MGPIO31B_H2F_B, I2C0_SDA_MGPIO30B_H2F_A, 
        I2C0_SDA_MGPIO30B_H2F_B, I2C1_SCL_MGPIO1A_H2F_A, 
        I2C1_SCL_MGPIO1A_H2F_B, I2C1_SDA_MGPIO0A_H2F_A, 
        I2C1_SDA_MGPIO0A_H2F_B, MDCF, MDOENF, MDOF, 
        MMUART0_CTS_MGPIO19B_H2F_A, MMUART0_CTS_MGPIO19B_H2F_B, 
        MMUART0_DCD_MGPIO22B_H2F_A, MMUART0_DCD_MGPIO22B_H2F_B, 
        MMUART0_DSR_MGPIO20B_H2F_A, MMUART0_DSR_MGPIO20B_H2F_B, 
        MMUART0_DTR_MGPIO18B_H2F_A, MMUART0_DTR_MGPIO18B_H2F_B, 
        MMUART0_RI_MGPIO21B_H2F_A, MMUART0_RI_MGPIO21B_H2F_B, 
        MMUART0_RTS_MGPIO17B_H2F_A, MMUART0_RTS_MGPIO17B_H2F_B, 
        MMUART0_RXD_MGPIO28B_H2F_A, MMUART0_RXD_MGPIO28B_H2F_B, 
        MMUART0_SCK_MGPIO29B_H2F_A, MMUART0_SCK_MGPIO29B_H2F_B, 
        MMUART0_TXD_MGPIO27B_H2F_A, MMUART0_TXD_MGPIO27B_H2F_B, 
        MMUART1_DTR_MGPIO12B_H2F_A, MMUART1_RTS_MGPIO11B_H2F_A, 
        MMUART1_RTS_MGPIO11B_H2F_B, MMUART1_RXD_MGPIO26B_H2F_A, 
        MMUART1_RXD_MGPIO26B_H2F_B, MMUART1_SCK_MGPIO25B_H2F_A, 
        MMUART1_SCK_MGPIO25B_H2F_B, MMUART1_TXD_MGPIO24B_H2F_A, 
        MMUART1_TXD_MGPIO24B_H2F_B, MPLL_LOCK, PER2_FABRIC_PENABLE, 
        PER2_FABRIC_PSEL, PER2_FABRIC_PWRITE, RTC_MATCH, SLEEPDEEP, 
        SLEEPHOLDACK, SLEEPING, SMBALERT_NO0, SMBALERT_NO1, SMBSUS_NO0, 
        SMBSUS_NO1, SPI0_CLK_OUT, SPI0_SDI_MGPIO5A_H2F_A, 
        SPI0_SDI_MGPIO5A_H2F_B, SPI0_SDO_MGPIO6A_H2F_A, 
        SPI0_SDO_MGPIO6A_H2F_B, SPI0_SS0_MGPIO7A_H2F_A, 
        SPI0_SS0_MGPIO7A_H2F_B, SPI0_SS1_MGPIO8A_H2F_A, 
        SPI0_SS1_MGPIO8A_H2F_B, SPI0_SS2_MGPIO9A_H2F_A, 
        SPI0_SS2_MGPIO9A_H2F_B, SPI0_SS3_MGPIO10A_H2F_A, 
        SPI0_SS3_MGPIO10A_H2F_B, SPI0_SS4_MGPIO19A_H2F_A, 
        SPI0_SS5_MGPIO20A_H2F_A, SPI0_SS6_MGPIO21A_H2F_A, 
        SPI0_SS7_MGPIO22A_H2F_A, SPI1_CLK_OUT, SPI1_SDI_MGPIO11A_H2F_A, 
        SPI1_SDI_MGPIO11A_H2F_B, SPI1_SDO_MGPIO12A_H2F_A, 
        SPI1_SDO_MGPIO12A_H2F_B, SPI1_SS0_MGPIO13A_H2F_A, 
        SPI1_SS0_MGPIO13A_H2F_B, SPI1_SS1_MGPIO14A_H2F_A, 
        SPI1_SS1_MGPIO14A_H2F_B, SPI1_SS2_MGPIO15A_H2F_A, 
        SPI1_SS2_MGPIO15A_H2F_B, SPI1_SS3_MGPIO16A_H2F_A, 
        SPI1_SS3_MGPIO16A_H2F_B, SPI1_SS4_MGPIO17A_H2F_A, 
        SPI1_SS5_MGPIO18A_H2F_A, SPI1_SS6_MGPIO23A_H2F_A, 
        SPI1_SS7_MGPIO24A_H2F_A, TRACECLK, TX_CLK, TXCTL_EN_RIF, TXEV, 
        WDOGTIMEOUT, F_ARREADY_HREADYOUT1, F_AWREADY_HREADYOUT0, 
        F_BVALID, F_RLAST, F_RVALID, F_WREADY, MDDR_FABRIC_PREADY, 
        MDDR_FABRIC_PSLVERR, VCC, GND, MDDR_DQS_0_PAD_Y, 
        MDDR_DQS_1_PAD_Y, CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT, MSS_ADLIB_INST_DRAM_CLK, 
        MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT, MMUART0_DCD_MGPIO22B_OUT, 
        MMUART0_DSR_MGPIO20B_OUT, MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT, 
        MMUART0_RI_MGPIO21B_OUT, MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT, 
        MMUART0_RXD_USBC_STP_MGPIO28B_OUT, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_OUT, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT, RGMII_MDC_RMII_MDC_OUT, 
        RGMII_RX_CLK_OUT, RGMII_TX_CLK_OUT, 
        RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT, 
        RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT, 
        SPI0_SDI_USBA_DIR_MGPIO5A_OUT, SPI0_SS1_USBA_DATA5_MGPIO8A_OUT, 
        SPI0_SS2_USBA_DATA6_MGPIO9A_OUT, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_OUT, SPI1_SDI_MGPIO11A_OUT, 
        SPI1_SS1_MGPIO14A_OUT, SPI1_SS2_MGPIO15A_OUT, 
        SPI1_SS3_MGPIO16A_OUT, SPI1_SS4_MGPIO17A_OUT, 
        SPI1_SS5_MGPIO18A_OUT, SPI1_SS6_MGPIO23A_OUT, 
        SPI1_SS7_MGPIO24A_OUT, USBC_XCLK_OUT, 
        CAN_RXBUS_USBA_DATA1_MGPIO3A_OE, 
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE, 
        CAN_TXBUS_USBA_DATA0_MGPIO2A_OE, 
        MMUART0_CTS_USBC_DATA7_MGPIO19B_OE, MMUART0_DCD_MGPIO22B_OE, 
        MMUART0_DSR_MGPIO20B_OE, MMUART0_DTR_USBC_DATA6_MGPIO18B_OE, 
        MMUART0_RI_MGPIO21B_OE, MMUART0_RTS_USBC_DATA5_MGPIO17B_OE, 
        MMUART0_RXD_USBC_STP_MGPIO28B_OE, 
        MMUART0_SCK_USBC_NXT_MGPIO29B_OE, 
        MMUART1_RXD_USBC_DATA3_MGPIO26B_OE, 
        MMUART1_SCK_USBC_DATA4_MGPIO25B_OE, 
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE, RGMII_MDC_RMII_MDC_OE, 
        RGMII_RX_CLK_OE, RGMII_TX_CLK_OE, 
        RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE, 
        RGMII_TXD0_RMII_TXD0_USBB_DIR_OE, SPI0_SDI_USBA_DIR_MGPIO5A_OE, 
        SPI0_SS1_USBA_DATA5_MGPIO8A_OE, SPI0_SS2_USBA_DATA6_MGPIO9A_OE, 
        SPI0_SS3_USBA_DATA7_MGPIO10A_OE, SPI1_SDI_MGPIO11A_OE, 
        SPI1_SS1_MGPIO14A_OE, SPI1_SS2_MGPIO15A_OE, 
        SPI1_SS3_MGPIO16A_OE, SPI1_SS4_MGPIO17A_OE, 
        SPI1_SS5_MGPIO18A_OE, SPI1_SS6_MGPIO23A_OE, 
        SPI1_SS7_MGPIO24A_OE, USBC_XCLK_OE;
    
    INBUF #( .IOSTD("") )  MMUART_0_RXD_PAD (.PAD(MMUART_0_RXD), .Y(
        MMUART_0_RXD_PAD_Y));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_ADDR_6_PAD (.D(
        DRAM_ADDR_net_0[6]), .PAD(MDDR_ADDR[6]));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_CAS_N_PAD (.D(
        MSS_ADLIB_INST_DRAM_CASN), .PAD(MDDR_CAS_N));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_RESET_N_PAD (.D(
        MSS_ADLIB_INST_DRAM_RSTN), .PAD(MDDR_RESET_N));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_ODT_PAD (.D(
        MSS_ADLIB_INST_DRAM_ODT), .PAD(MDDR_ODT));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_ADDR_11_PAD (.D(
        DRAM_ADDR_net_0[11]), .PAD(MDDR_ADDR[11]));
    TRIBUFF #( .IOSTD("") )  MMUART_1_TXD_PAD (.D(
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT), .E(
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OE), .PAD(
        MMUART_1_TXD));
    BIBUF #( .IOSTD("SSTL18I") )  MDDR_DQ_10_PAD (.PAD(MDDR_DQ[10]), 
        .D(DRAM_DQ_OUT_net_0[10]), .E(DRAM_DQ_OE_net_0[10]), .Y(
        MDDR_DQ_10_PAD_Y));
    INBUF #( .IOSTD("") )  USB_ULPI_XCLK_PAD (.PAD(USB_ULPI_XCLK), .Y(
        USB_ULPI_XCLK_PAD_Y));
    BIBUF #( .IOSTD("SSTL18I") )  MDDR_DQ_1_PAD (.PAD(MDDR_DQ[1]), .D(
        DRAM_DQ_OUT_net_0[1]), .E(DRAM_DQ_OE_net_0[1]), .Y(
        MDDR_DQ_1_PAD_Y));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_ADDR_7_PAD (.D(
        DRAM_ADDR_net_0[7]), .PAD(MDDR_ADDR[7]));
    BIBUF #( .IOSTD("SSTL18I") )  MDDR_DQ_11_PAD (.PAD(MDDR_DQ[11]), 
        .D(DRAM_DQ_OUT_net_0[11]), .E(DRAM_DQ_OE_net_0[11]), .Y(
        MDDR_DQ_11_PAD_Y));
    INBUF #( .IOSTD("") )  USB_ULPI_DIR_PAD (.PAD(USB_ULPI_DIR), .Y(
        USB_ULPI_DIR_PAD_Y));
    BIBUF #( .IOSTD("SSTL18I") )  MDDR_DQ_9_PAD (.PAD(MDDR_DQ[9]), .D(
        DRAM_DQ_OUT_net_0[9]), .E(DRAM_DQ_OE_net_0[9]), .Y(
        MDDR_DQ_9_PAD_Y));
    BIBUF #( .IOSTD("SSTL18I") )  MDDR_DQ_3_PAD (.PAD(MDDR_DQ[3]), .D(
        DRAM_DQ_OUT_net_0[3]), .E(DRAM_DQ_OE_net_0[3]), .Y(
        MDDR_DQ_3_PAD_Y));
    BIBUF #( .IOSTD("SSTL18I") )  MDDR_DQ_0_PAD (.PAD(MDDR_DQ[0]), .D(
        DRAM_DQ_OUT_net_0[0]), .E(DRAM_DQ_OE_net_0[0]), .Y(
        MDDR_DQ_0_PAD_Y));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_ADDR_12_PAD (.D(
        DRAM_ADDR_net_0[12]), .PAD(MDDR_ADDR[12]));
    BIBUF #( .IOSTD("") )  USB_ULPI_DATA_2_PAD (.PAD(USB_ULPI_DATA[2]), 
        .D(MSS_ADLIB_INST_RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT), .E(
        MSS_ADLIB_INST_RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE), .Y(
        USB_ULPI_DATA_2_PAD_Y));
    BIBUF #( .IOSTD("") )  SPI_1_SS0_PAD (.PAD(SPI_1_SS0), .D(
        MSS_ADLIB_INST_SPI1_SS0_MGPIO13A_OUT), .E(
        MSS_ADLIB_INST_SPI1_SS0_MGPIO13A_OE), .Y(SPI_1_SS0_PAD_Y));
    BIBUF #( .IOSTD("SSTL18I") )  MDDR_DQ_2_PAD (.PAD(MDDR_DQ[2]), .D(
        DRAM_DQ_OUT_net_0[2]), .E(DRAM_DQ_OE_net_0[2]), .Y(
        MDDR_DQ_2_PAD_Y));
    BIBUF #( .IOSTD("SSTL18I") )  MDDR_DQ_12_PAD (.PAD(MDDR_DQ[12]), 
        .D(DRAM_DQ_OUT_net_0[12]), .E(DRAM_DQ_OE_net_0[12]), .Y(
        MDDR_DQ_12_PAD_Y));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_CKE_PAD (.D(
        MSS_ADLIB_INST_DRAM_CKE), .PAD(MDDR_CKE));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_ADDR_2_PAD (.D(
        DRAM_ADDR_net_0[2]), .PAD(MDDR_ADDR[2]));
    TRIBUFF #( .IOSTD("") )  MMUART_0_TXD_PAD (.D(
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OUT), .E(
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OE), .PAD(
        MMUART_0_TXD));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_ADDR_13_PAD (.D(
        DRAM_ADDR_net_0[13]), .PAD(MDDR_ADDR[13]));
    BIBUF #( .IOSTD("") )  I2C_1_SDA_PAD (.PAD(I2C_1_SDA), .D(
        MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OUT), .E(
        MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OE), .Y(
        I2C_1_SDA_PAD_Y));
    BIBUF #( .IOSTD("") )  USB_ULPI_DATA_0_PAD (.PAD(USB_ULPI_DATA[0]), 
        .D(MSS_ADLIB_INST_RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT), .E(
        MSS_ADLIB_INST_RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE), .Y(
        USB_ULPI_DATA_0_PAD_Y));
    BIBUF #( .IOSTD("") )  I2C_1_SCL_PAD (.PAD(I2C_1_SCL), .D(
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OUT), .E(
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OE), .Y(
        I2C_1_SCL_PAD_Y));
    BIBUF #( .IOSTD("") )  USB_ULPI_DATA_7_PAD (.PAD(USB_ULPI_DATA[7]), 
        .D(MSS_ADLIB_INST_RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT), .E(
        MSS_ADLIB_INST_RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE), .Y(
        USB_ULPI_DATA_7_PAD_Y));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_ADDR_5_PAD (.D(
        DRAM_ADDR_net_0[5]), .PAD(MDDR_ADDR[5]));
    TRIBUFF #( .IOSTD("") )  SPI_1_DO_PAD (.D(
        MSS_ADLIB_INST_SPI1_SDO_MGPIO12A_OUT), .E(
        MSS_ADLIB_INST_SPI1_SDO_MGPIO12A_OE), .PAD(SPI_1_DO));
    BIBUF #( .IOSTD("SSTL18I") )  MDDR_DM_RDQS_1_PAD (.PAD(
        MDDR_DM_RDQS[1]), .D(DRAM_DM_RDQS_OUT_net_0[1]), .E(
        DM_OE_net_0[1]), .Y(MDDR_DM_RDQS_1_PAD_Y));
    TRIBUFF #( .IOSTD("") )  SPI_0_DO_PAD (.D(
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OUT), .E(
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OE), .PAD(SPI_0_DO));
    BIBUF_DIFF #( .IOSTD("SSTL18I") )  MDDR_DQS_0_PAD (.D(
        DRAM_DQS_OUT_net_0[0]), .E(DRAM_DQS_OE_net_0[0]), .PADP(
        MDDR_DQS[0]), .PADN(MDDR_DQS_N[0]), .Y(MDDR_DQS_0_PAD_Y));
    BIBUF_DIFF #( .IOSTD("SSTL18I") )  MDDR_DQS_1_PAD (.D(
        DRAM_DQS_OUT_net_0[1]), .E(DRAM_DQS_OE_net_0[1]), .PADP(
        MDDR_DQS[1]), .PADN(MDDR_DQS_N[1]), .Y(MDDR_DQS_1_PAD_Y));
    BIBUF #( .IOSTD("SSTL18I") )  MDDR_DQ_15_PAD (.PAD(MDDR_DQ[15]), 
        .D(DRAM_DQ_OUT_net_0[15]), .E(DRAM_DQ_OE_net_0[15]), .Y(
        MDDR_DQ_15_PAD_Y));
    BIBUF #( .IOSTD("SSTL18I") )  MDDR_DM_RDQS_0_PAD (.PAD(
        MDDR_DM_RDQS[0]), .D(DRAM_DM_RDQS_OUT_net_0[0]), .E(
        DM_OE_net_0[0]), .Y(MDDR_DM_RDQS_0_PAD_Y));
    INBUF #( .IOSTD("") )  SPI_1_DI_PAD (.PAD(SPI_1_DI), .Y(
        SPI_1_DI_PAD_Y));
    BIBUF #( .IOSTD("") )  I2C_0_SCL_PAD (.PAD(I2C_0_SCL), .D(
        MSS_ADLIB_INST_I2C0_SCL_USBC_DATA1_MGPIO31B_OUT), .E(
        MSS_ADLIB_INST_I2C0_SCL_USBC_DATA1_MGPIO31B_OE), .Y(
        I2C_0_SCL_PAD_Y));
    INBUF #( .IOSTD("") )  SPI_0_DI_PAD (.PAD(SPI_0_DI), .Y(
        SPI_0_DI_PAD_Y));
    BIBUF #( .IOSTD("SSTL18I") )  MDDR_DQ_8_PAD (.PAD(MDDR_DQ[8]), .D(
        DRAM_DQ_OUT_net_0[8]), .E(DRAM_DQ_OE_net_0[8]), .Y(
        MDDR_DQ_8_PAD_Y));
    TRIBUFF #( .IOSTD("") )  USB_ULPI_STP_PAD (.D(
        MSS_ADLIB_INST_RGMII_TXD1_RMII_TXD1_USBB_STP_OUT), .E(
        MSS_ADLIB_INST_RGMII_TXD1_RMII_TXD1_USBB_STP_OE), .PAD(
        USB_ULPI_STP));
    BIBUF #( .IOSTD("") )  USB_ULPI_DATA_4_PAD (.PAD(USB_ULPI_DATA[4]), 
        .D(MSS_ADLIB_INST_RGMII_RXD3_USBB_DATA4_OUT), .E(
        MSS_ADLIB_INST_RGMII_RXD3_USBB_DATA4_OE), .Y(
        USB_ULPI_DATA_4_PAD_Y));
    BIBUF #( .IOSTD("") )  USB_ULPI_DATA_3_PAD (.PAD(USB_ULPI_DATA[3]), 
        .D(MSS_ADLIB_INST_RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT), .E(
        MSS_ADLIB_INST_RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE), .Y(
        USB_ULPI_DATA_3_PAD_Y));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_ADDR_9_PAD (.D(
        DRAM_ADDR_net_0[9]), .PAD(MDDR_ADDR[9]));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_BA_2_PAD (.D(DRAM_BA_net_0[2]), 
        .PAD(MDDR_BA[2]));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_ADDR_14_PAD (.D(
        DRAM_ADDR_net_0[14]), .PAD(MDDR_ADDR[14]));
    MSS_010 #( .INIT(1438'h0000040100361200000000000000003610008000000000000000000000000000000000001203610000000000000000000120361000000000100520481204812048120D8120D8120F00000000F000000000000000000000000000000007FFFFFFFB000001007C37F00020200E09280F00183FFFFE400000000002150000000000E11C0000007E4800010842108421000001FE34001FF8000000400000000020091007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
        , .ACT_UBITS(56'b11111111111111111111111111111111111111111111111111111111)
        , .MEMORYFILE("ENVM_init.mem"), .RTC_MAIN_XTL_FREQ(0.000000), .RTC_MAIN_XTL_MODE("")
        , .DDR_CLK_FREQ(200.000000) )  MSS_ADLIB_INST (
        .CAN_RXBUS_MGPIO3A_H2F_A(CAN_RXBUS_MGPIO3A_H2F_A), 
        .CAN_RXBUS_MGPIO3A_H2F_B(CAN_RXBUS_MGPIO3A_H2F_B), 
        .CAN_TX_EBL_MGPIO4A_H2F_A(CAN_TX_EBL_MGPIO4A_H2F_A), 
        .CAN_TX_EBL_MGPIO4A_H2F_B(CAN_TX_EBL_MGPIO4A_H2F_B), 
        .CAN_TXBUS_MGPIO2A_H2F_A(CAN_TXBUS_MGPIO2A_H2F_A), 
        .CAN_TXBUS_MGPIO2A_H2F_B(CAN_TXBUS_MGPIO2A_H2F_B), 
        .CLK_CONFIG_APB(CLK_CONFIG_APB), .COMMS_INT(COMMS_INT), 
        .CONFIG_PRESET_N(CONFIG_PRESET_N), .EDAC_ERROR({EDAC_ERROR[7], 
        EDAC_ERROR[6], EDAC_ERROR[5], EDAC_ERROR[4], EDAC_ERROR[3], 
        EDAC_ERROR[2], EDAC_ERROR[1], EDAC_ERROR[0]}), .F_FM0_RDATA({
        F_FM0_RDATA[31], F_FM0_RDATA[30], F_FM0_RDATA[29], 
        F_FM0_RDATA[28], F_FM0_RDATA[27], F_FM0_RDATA[26], 
        F_FM0_RDATA[25], F_FM0_RDATA[24], F_FM0_RDATA[23], 
        F_FM0_RDATA[22], F_FM0_RDATA[21], F_FM0_RDATA[20], 
        F_FM0_RDATA[19], F_FM0_RDATA[18], F_FM0_RDATA[17], 
        F_FM0_RDATA[16], F_FM0_RDATA[15], F_FM0_RDATA[14], 
        F_FM0_RDATA[13], F_FM0_RDATA[12], F_FM0_RDATA[11], 
        F_FM0_RDATA[10], F_FM0_RDATA[9], F_FM0_RDATA[8], 
        F_FM0_RDATA[7], F_FM0_RDATA[6], F_FM0_RDATA[5], F_FM0_RDATA[4], 
        F_FM0_RDATA[3], F_FM0_RDATA[2], F_FM0_RDATA[1], F_FM0_RDATA[0]})
        , .F_FM0_READYOUT(F_FM0_READYOUT), .F_FM0_RESP(F_FM0_RESP), 
        .F_HM0_ADDR({F_HM0_ADDR[31], F_HM0_ADDR[30], F_HM0_ADDR[29], 
        F_HM0_ADDR[28], F_HM0_ADDR[27], F_HM0_ADDR[26], F_HM0_ADDR[25], 
        F_HM0_ADDR[24], F_HM0_ADDR[23], F_HM0_ADDR[22], F_HM0_ADDR[21], 
        F_HM0_ADDR[20], F_HM0_ADDR[19], F_HM0_ADDR[18], F_HM0_ADDR[17], 
        F_HM0_ADDR[16], F_HM0_ADDR[15], F_HM0_ADDR[14], F_HM0_ADDR[13], 
        F_HM0_ADDR[12], F_HM0_ADDR[11], F_HM0_ADDR[10], F_HM0_ADDR[9], 
        F_HM0_ADDR[8], F_HM0_ADDR[7], F_HM0_ADDR[6], F_HM0_ADDR[5], 
        F_HM0_ADDR[4], F_HM0_ADDR[3], F_HM0_ADDR[2], F_HM0_ADDR[1], 
        F_HM0_ADDR[0]}), .F_HM0_ENABLE(F_HM0_ENABLE), .F_HM0_SEL(
        F_HM0_SEL), .F_HM0_SIZE({F_HM0_SIZE[1], F_HM0_SIZE[0]}), 
        .F_HM0_TRANS1(F_HM0_TRANS1), .F_HM0_WDATA({F_HM0_WDATA[31], 
        F_HM0_WDATA[30], F_HM0_WDATA[29], F_HM0_WDATA[28], 
        F_HM0_WDATA[27], F_HM0_WDATA[26], F_HM0_WDATA[25], 
        F_HM0_WDATA[24], F_HM0_WDATA[23], F_HM0_WDATA[22], 
        F_HM0_WDATA[21], F_HM0_WDATA[20], F_HM0_WDATA[19], 
        F_HM0_WDATA[18], F_HM0_WDATA[17], F_HM0_WDATA[16], 
        F_HM0_WDATA[15], F_HM0_WDATA[14], F_HM0_WDATA[13], 
        F_HM0_WDATA[12], F_HM0_WDATA[11], F_HM0_WDATA[10], 
        F_HM0_WDATA[9], F_HM0_WDATA[8], F_HM0_WDATA[7], F_HM0_WDATA[6], 
        F_HM0_WDATA[5], F_HM0_WDATA[4], F_HM0_WDATA[3], F_HM0_WDATA[2], 
        F_HM0_WDATA[1], F_HM0_WDATA[0]}), .F_HM0_WRITE(F_HM0_WRITE), 
        .FAB_CHRGVBUS(FAB_CHRGVBUS), .FAB_DISCHRGVBUS(FAB_DISCHRGVBUS), 
        .FAB_DMPULLDOWN(FAB_DMPULLDOWN), .FAB_DPPULLDOWN(
        FAB_DPPULLDOWN), .FAB_DRVVBUS(FAB_DRVVBUS), .FAB_IDPULLUP(
        FAB_IDPULLUP), .FAB_OPMODE({FAB_OPMODE[1], FAB_OPMODE[0]}), 
        .FAB_SUSPENDM(FAB_SUSPENDM), .FAB_TERMSEL(FAB_TERMSEL), 
        .FAB_TXVALID(FAB_TXVALID), .FAB_VCONTROL({FAB_VCONTROL[3], 
        FAB_VCONTROL[2], FAB_VCONTROL[1], FAB_VCONTROL[0]}), 
        .FAB_VCONTROLLOADM(FAB_VCONTROLLOADM), .FAB_XCVRSEL({
        FAB_XCVRSEL[1], FAB_XCVRSEL[0]}), .FAB_XDATAOUT({
        FAB_XDATAOUT[7], FAB_XDATAOUT[6], FAB_XDATAOUT[5], 
        FAB_XDATAOUT[4], FAB_XDATAOUT[3], FAB_XDATAOUT[2], 
        FAB_XDATAOUT[1], FAB_XDATAOUT[0]}), .FACC_GLMUX_SEL(
        FACC_GLMUX_SEL), .FIC32_0_MASTER({FIC32_0_MASTER[1], 
        FIC32_0_MASTER[0]}), .FIC32_1_MASTER({FIC32_1_MASTER[1], 
        FIC32_1_MASTER[0]}), .FPGA_RESET_N(FPGA_RESET_N), .GTX_CLK(
        GTX_CLK), .H2F_INTERRUPT({H2F_INTERRUPT[15], H2F_INTERRUPT[14], 
        H2F_INTERRUPT[13], H2F_INTERRUPT[12], H2F_INTERRUPT[11], 
        H2F_INTERRUPT[10], H2F_INTERRUPT[9], H2F_INTERRUPT[8], 
        H2F_INTERRUPT[7], H2F_INTERRUPT[6], H2F_INTERRUPT[5], 
        H2F_INTERRUPT[4], H2F_INTERRUPT[3], H2F_INTERRUPT[2], 
        H2F_INTERRUPT[1], H2F_INTERRUPT[0]}), .H2F_NMI(H2F_NMI), 
        .H2FCALIB(H2FCALIB), .I2C0_SCL_MGPIO31B_H2F_A(
        I2C0_SCL_MGPIO31B_H2F_A), .I2C0_SCL_MGPIO31B_H2F_B(
        I2C0_SCL_MGPIO31B_H2F_B), .I2C0_SDA_MGPIO30B_H2F_A(
        I2C0_SDA_MGPIO30B_H2F_A), .I2C0_SDA_MGPIO30B_H2F_B(
        I2C0_SDA_MGPIO30B_H2F_B), .I2C1_SCL_MGPIO1A_H2F_A(
        I2C1_SCL_MGPIO1A_H2F_A), .I2C1_SCL_MGPIO1A_H2F_B(
        I2C1_SCL_MGPIO1A_H2F_B), .I2C1_SDA_MGPIO0A_H2F_A(
        I2C1_SDA_MGPIO0A_H2F_A), .I2C1_SDA_MGPIO0A_H2F_B(
        I2C1_SDA_MGPIO0A_H2F_B), .MDCF(MDCF), .MDOENF(MDOENF), .MDOF(
        MDOF), .MMUART0_CTS_MGPIO19B_H2F_A(MMUART0_CTS_MGPIO19B_H2F_A), 
        .MMUART0_CTS_MGPIO19B_H2F_B(MMUART0_CTS_MGPIO19B_H2F_B), 
        .MMUART0_DCD_MGPIO22B_H2F_A(MMUART0_DCD_MGPIO22B_H2F_A), 
        .MMUART0_DCD_MGPIO22B_H2F_B(MMUART0_DCD_MGPIO22B_H2F_B), 
        .MMUART0_DSR_MGPIO20B_H2F_A(MMUART0_DSR_MGPIO20B_H2F_A), 
        .MMUART0_DSR_MGPIO20B_H2F_B(MMUART0_DSR_MGPIO20B_H2F_B), 
        .MMUART0_DTR_MGPIO18B_H2F_A(MMUART0_DTR_MGPIO18B_H2F_A), 
        .MMUART0_DTR_MGPIO18B_H2F_B(MMUART0_DTR_MGPIO18B_H2F_B), 
        .MMUART0_RI_MGPIO21B_H2F_A(MMUART0_RI_MGPIO21B_H2F_A), 
        .MMUART0_RI_MGPIO21B_H2F_B(MMUART0_RI_MGPIO21B_H2F_B), 
        .MMUART0_RTS_MGPIO17B_H2F_A(MMUART0_RTS_MGPIO17B_H2F_A), 
        .MMUART0_RTS_MGPIO17B_H2F_B(MMUART0_RTS_MGPIO17B_H2F_B), 
        .MMUART0_RXD_MGPIO28B_H2F_A(MMUART0_RXD_MGPIO28B_H2F_A), 
        .MMUART0_RXD_MGPIO28B_H2F_B(MMUART0_RXD_MGPIO28B_H2F_B), 
        .MMUART0_SCK_MGPIO29B_H2F_A(MMUART0_SCK_MGPIO29B_H2F_A), 
        .MMUART0_SCK_MGPIO29B_H2F_B(MMUART0_SCK_MGPIO29B_H2F_B), 
        .MMUART0_TXD_MGPIO27B_H2F_A(MMUART0_TXD_MGPIO27B_H2F_A), 
        .MMUART0_TXD_MGPIO27B_H2F_B(MMUART0_TXD_MGPIO27B_H2F_B), 
        .MMUART1_DTR_MGPIO12B_H2F_A(MMUART1_DTR_MGPIO12B_H2F_A), 
        .MMUART1_RTS_MGPIO11B_H2F_A(MMUART1_RTS_MGPIO11B_H2F_A), 
        .MMUART1_RTS_MGPIO11B_H2F_B(MMUART1_RTS_MGPIO11B_H2F_B), 
        .MMUART1_RXD_MGPIO26B_H2F_A(MMUART1_RXD_MGPIO26B_H2F_A), 
        .MMUART1_RXD_MGPIO26B_H2F_B(MMUART1_RXD_MGPIO26B_H2F_B), 
        .MMUART1_SCK_MGPIO25B_H2F_A(MMUART1_SCK_MGPIO25B_H2F_A), 
        .MMUART1_SCK_MGPIO25B_H2F_B(MMUART1_SCK_MGPIO25B_H2F_B), 
        .MMUART1_TXD_MGPIO24B_H2F_A(MMUART1_TXD_MGPIO24B_H2F_A), 
        .MMUART1_TXD_MGPIO24B_H2F_B(MMUART1_TXD_MGPIO24B_H2F_B), 
        .MPLL_LOCK(MPLL_LOCK), .PER2_FABRIC_PADDR({
        PER2_FABRIC_PADDR[15], PER2_FABRIC_PADDR[14], 
        PER2_FABRIC_PADDR[13], PER2_FABRIC_PADDR[12], 
        PER2_FABRIC_PADDR[11], PER2_FABRIC_PADDR[10], 
        PER2_FABRIC_PADDR[9], PER2_FABRIC_PADDR[8], 
        PER2_FABRIC_PADDR[7], PER2_FABRIC_PADDR[6], 
        PER2_FABRIC_PADDR[5], PER2_FABRIC_PADDR[4], 
        PER2_FABRIC_PADDR[3], PER2_FABRIC_PADDR[2]}), 
        .PER2_FABRIC_PENABLE(PER2_FABRIC_PENABLE), .PER2_FABRIC_PSEL(
        PER2_FABRIC_PSEL), .PER2_FABRIC_PWDATA({PER2_FABRIC_PWDATA[31], 
        PER2_FABRIC_PWDATA[30], PER2_FABRIC_PWDATA[29], 
        PER2_FABRIC_PWDATA[28], PER2_FABRIC_PWDATA[27], 
        PER2_FABRIC_PWDATA[26], PER2_FABRIC_PWDATA[25], 
        PER2_FABRIC_PWDATA[24], PER2_FABRIC_PWDATA[23], 
        PER2_FABRIC_PWDATA[22], PER2_FABRIC_PWDATA[21], 
        PER2_FABRIC_PWDATA[20], PER2_FABRIC_PWDATA[19], 
        PER2_FABRIC_PWDATA[18], PER2_FABRIC_PWDATA[17], 
        PER2_FABRIC_PWDATA[16], PER2_FABRIC_PWDATA[15], 
        PER2_FABRIC_PWDATA[14], PER2_FABRIC_PWDATA[13], 
        PER2_FABRIC_PWDATA[12], PER2_FABRIC_PWDATA[11], 
        PER2_FABRIC_PWDATA[10], PER2_FABRIC_PWDATA[9], 
        PER2_FABRIC_PWDATA[8], PER2_FABRIC_PWDATA[7], 
        PER2_FABRIC_PWDATA[6], PER2_FABRIC_PWDATA[5], 
        PER2_FABRIC_PWDATA[4], PER2_FABRIC_PWDATA[3], 
        PER2_FABRIC_PWDATA[2], PER2_FABRIC_PWDATA[1], 
        PER2_FABRIC_PWDATA[0]}), .PER2_FABRIC_PWRITE(
        PER2_FABRIC_PWRITE), .RTC_MATCH(RTC_MATCH), .SLEEPDEEP(
        SLEEPDEEP), .SLEEPHOLDACK(SLEEPHOLDACK), .SLEEPING(SLEEPING), 
        .SMBALERT_NO0(SMBALERT_NO0), .SMBALERT_NO1(SMBALERT_NO1), 
        .SMBSUS_NO0(SMBSUS_NO0), .SMBSUS_NO1(SMBSUS_NO1), 
        .SPI0_CLK_OUT(SPI0_CLK_OUT), .SPI0_SDI_MGPIO5A_H2F_A(
        SPI0_SDI_MGPIO5A_H2F_A), .SPI0_SDI_MGPIO5A_H2F_B(
        SPI0_SDI_MGPIO5A_H2F_B), .SPI0_SDO_MGPIO6A_H2F_A(
        SPI0_SDO_MGPIO6A_H2F_A), .SPI0_SDO_MGPIO6A_H2F_B(
        SPI0_SDO_MGPIO6A_H2F_B), .SPI0_SS0_MGPIO7A_H2F_A(
        SPI0_SS0_MGPIO7A_H2F_A), .SPI0_SS0_MGPIO7A_H2F_B(
        SPI0_SS0_MGPIO7A_H2F_B), .SPI0_SS1_MGPIO8A_H2F_A(
        SPI0_SS1_MGPIO8A_H2F_A), .SPI0_SS1_MGPIO8A_H2F_B(
        SPI0_SS1_MGPIO8A_H2F_B), .SPI0_SS2_MGPIO9A_H2F_A(
        SPI0_SS2_MGPIO9A_H2F_A), .SPI0_SS2_MGPIO9A_H2F_B(
        SPI0_SS2_MGPIO9A_H2F_B), .SPI0_SS3_MGPIO10A_H2F_A(
        SPI0_SS3_MGPIO10A_H2F_A), .SPI0_SS3_MGPIO10A_H2F_B(
        SPI0_SS3_MGPIO10A_H2F_B), .SPI0_SS4_MGPIO19A_H2F_A(
        SPI0_SS4_MGPIO19A_H2F_A), .SPI0_SS5_MGPIO20A_H2F_A(
        SPI0_SS5_MGPIO20A_H2F_A), .SPI0_SS6_MGPIO21A_H2F_A(
        SPI0_SS6_MGPIO21A_H2F_A), .SPI0_SS7_MGPIO22A_H2F_A(
        SPI0_SS7_MGPIO22A_H2F_A), .SPI1_CLK_OUT(SPI1_CLK_OUT), 
        .SPI1_SDI_MGPIO11A_H2F_A(SPI1_SDI_MGPIO11A_H2F_A), 
        .SPI1_SDI_MGPIO11A_H2F_B(SPI1_SDI_MGPIO11A_H2F_B), 
        .SPI1_SDO_MGPIO12A_H2F_A(SPI1_SDO_MGPIO12A_H2F_A), 
        .SPI1_SDO_MGPIO12A_H2F_B(SPI1_SDO_MGPIO12A_H2F_B), 
        .SPI1_SS0_MGPIO13A_H2F_A(SPI1_SS0_MGPIO13A_H2F_A), 
        .SPI1_SS0_MGPIO13A_H2F_B(SPI1_SS0_MGPIO13A_H2F_B), 
        .SPI1_SS1_MGPIO14A_H2F_A(SPI1_SS1_MGPIO14A_H2F_A), 
        .SPI1_SS1_MGPIO14A_H2F_B(SPI1_SS1_MGPIO14A_H2F_B), 
        .SPI1_SS2_MGPIO15A_H2F_A(SPI1_SS2_MGPIO15A_H2F_A), 
        .SPI1_SS2_MGPIO15A_H2F_B(SPI1_SS2_MGPIO15A_H2F_B), 
        .SPI1_SS3_MGPIO16A_H2F_A(SPI1_SS3_MGPIO16A_H2F_A), 
        .SPI1_SS3_MGPIO16A_H2F_B(SPI1_SS3_MGPIO16A_H2F_B), 
        .SPI1_SS4_MGPIO17A_H2F_A(SPI1_SS4_MGPIO17A_H2F_A), 
        .SPI1_SS5_MGPIO18A_H2F_A(SPI1_SS5_MGPIO18A_H2F_A), 
        .SPI1_SS6_MGPIO23A_H2F_A(SPI1_SS6_MGPIO23A_H2F_A), 
        .SPI1_SS7_MGPIO24A_H2F_A(SPI1_SS7_MGPIO24A_H2F_A), .TCGF({
        TCGF[9], TCGF[8], TCGF[7], TCGF[6], TCGF[5], TCGF[4], TCGF[3], 
        TCGF[2], TCGF[1], TCGF[0]}), .TRACECLK(TRACECLK), .TRACEDATA({
        TRACEDATA[3], TRACEDATA[2], TRACEDATA[1], TRACEDATA[0]}), 
        .TX_CLK(TX_CLK), .TX_ENF(MAC_MII_TX_EN), .TX_ERRF(
        MAC_MII_TX_ER), .TXCTL_EN_RIF(TXCTL_EN_RIF), .TXD_RIF({
        TXD_RIF[3], TXD_RIF[2], TXD_RIF[1], TXD_RIF[0]}), .TXDF({
        TXDF_net_0[7], TXDF_net_0[6], TXDF_net_0[5], TXDF_net_0[4], 
        MAC_MII_TXD[3], MAC_MII_TXD[2], MAC_MII_TXD[1], MAC_MII_TXD[0]})
        , .TXEV(TXEV), .WDOGTIMEOUT(WDOGTIMEOUT), 
        .F_ARREADY_HREADYOUT1(F_ARREADY_HREADYOUT1), 
        .F_AWREADY_HREADYOUT0(F_AWREADY_HREADYOUT0), .F_BID({F_BID[3], 
        F_BID[2], F_BID[1], F_BID[0]}), .F_BRESP_HRESP0({
        F_BRESP_HRESP0[1], F_BRESP_HRESP0[0]}), .F_BVALID(F_BVALID), 
        .F_RDATA_HRDATA01({F_RDATA_HRDATA01[63], F_RDATA_HRDATA01[62], 
        F_RDATA_HRDATA01[61], F_RDATA_HRDATA01[60], 
        F_RDATA_HRDATA01[59], F_RDATA_HRDATA01[58], 
        F_RDATA_HRDATA01[57], F_RDATA_HRDATA01[56], 
        F_RDATA_HRDATA01[55], F_RDATA_HRDATA01[54], 
        F_RDATA_HRDATA01[53], F_RDATA_HRDATA01[52], 
        F_RDATA_HRDATA01[51], F_RDATA_HRDATA01[50], 
        F_RDATA_HRDATA01[49], F_RDATA_HRDATA01[48], 
        F_RDATA_HRDATA01[47], F_RDATA_HRDATA01[46], 
        F_RDATA_HRDATA01[45], F_RDATA_HRDATA01[44], 
        F_RDATA_HRDATA01[43], F_RDATA_HRDATA01[42], 
        F_RDATA_HRDATA01[41], F_RDATA_HRDATA01[40], 
        F_RDATA_HRDATA01[39], F_RDATA_HRDATA01[38], 
        F_RDATA_HRDATA01[37], F_RDATA_HRDATA01[36], 
        F_RDATA_HRDATA01[35], F_RDATA_HRDATA01[34], 
        F_RDATA_HRDATA01[33], F_RDATA_HRDATA01[32], 
        F_RDATA_HRDATA01[31], F_RDATA_HRDATA01[30], 
        F_RDATA_HRDATA01[29], F_RDATA_HRDATA01[28], 
        F_RDATA_HRDATA01[27], F_RDATA_HRDATA01[26], 
        F_RDATA_HRDATA01[25], F_RDATA_HRDATA01[24], 
        F_RDATA_HRDATA01[23], F_RDATA_HRDATA01[22], 
        F_RDATA_HRDATA01[21], F_RDATA_HRDATA01[20], 
        F_RDATA_HRDATA01[19], F_RDATA_HRDATA01[18], 
        F_RDATA_HRDATA01[17], F_RDATA_HRDATA01[16], 
        F_RDATA_HRDATA01[15], F_RDATA_HRDATA01[14], 
        F_RDATA_HRDATA01[13], F_RDATA_HRDATA01[12], 
        F_RDATA_HRDATA01[11], F_RDATA_HRDATA01[10], 
        F_RDATA_HRDATA01[9], F_RDATA_HRDATA01[8], F_RDATA_HRDATA01[7], 
        F_RDATA_HRDATA01[6], F_RDATA_HRDATA01[5], F_RDATA_HRDATA01[4], 
        F_RDATA_HRDATA01[3], F_RDATA_HRDATA01[2], F_RDATA_HRDATA01[1], 
        F_RDATA_HRDATA01[0]}), .F_RID({F_RID[3], F_RID[2], F_RID[1], 
        F_RID[0]}), .F_RLAST(F_RLAST), .F_RRESP_HRESP1({
        F_RRESP_HRESP1[1], F_RRESP_HRESP1[0]}), .F_RVALID(F_RVALID), 
        .F_WREADY(F_WREADY), .MDDR_FABRIC_PRDATA({
        MDDR_FABRIC_PRDATA[15], MDDR_FABRIC_PRDATA[14], 
        MDDR_FABRIC_PRDATA[13], MDDR_FABRIC_PRDATA[12], 
        MDDR_FABRIC_PRDATA[11], MDDR_FABRIC_PRDATA[10], 
        MDDR_FABRIC_PRDATA[9], MDDR_FABRIC_PRDATA[8], 
        MDDR_FABRIC_PRDATA[7], MDDR_FABRIC_PRDATA[6], 
        MDDR_FABRIC_PRDATA[5], MDDR_FABRIC_PRDATA[4], 
        MDDR_FABRIC_PRDATA[3], MDDR_FABRIC_PRDATA[2], 
        MDDR_FABRIC_PRDATA[1], MDDR_FABRIC_PRDATA[0]}), 
        .MDDR_FABRIC_PREADY(MDDR_FABRIC_PREADY), .MDDR_FABRIC_PSLVERR(
        MDDR_FABRIC_PSLVERR), .CAN_RXBUS_F2H_SCP(VCC), 
        .CAN_TX_EBL_F2H_SCP(VCC), .CAN_TXBUS_F2H_SCP(VCC), .COLF(
        MAC_MII_COL), .CRSF(MAC_MII_CRS), .F2_DMAREADY({VCC, VCC}), 
        .F2H_INTERRUPT({GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND}), .F2HCALIB(VCC), 
        .F_DMAREADY({VCC, VCC}), .F_FM0_ADDR({GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND}), .F_FM0_ENABLE(GND), .F_FM0_MASTLOCK(GND), 
        .F_FM0_READY(VCC), .F_FM0_SEL(GND), .F_FM0_SIZE({GND, GND}), 
        .F_FM0_TRANS1(GND), .F_FM0_WDATA({GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND}), .F_FM0_WRITE(GND), .F_HM0_RDATA({GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND}), .F_HM0_READY(VCC), .F_HM0_RESP(GND), 
        .FAB_AVALID(VCC), .FAB_HOSTDISCON(VCC), .FAB_IDDIG(VCC), 
        .FAB_LINESTATE({VCC, VCC}), .FAB_M3_RESET_N(VCC), 
        .FAB_PLL_LOCK(VCC), .FAB_RXACTIVE(VCC), .FAB_RXERROR(VCC), 
        .FAB_RXVALID(VCC), .FAB_RXVALIDH(GND), .FAB_SESSEND(VCC), 
        .FAB_TXREADY(VCC), .FAB_VBUSVALID(VCC), .FAB_VSTATUS({VCC, VCC, 
        VCC, VCC, VCC, VCC, VCC, VCC}), .FAB_XDATAIN({VCC, VCC, VCC, 
        VCC, VCC, VCC, VCC, VCC}), .GTX_CLKPF(VCC), .I2C0_BCLK(VCC), 
        .I2C0_SCL_F2H_SCP(VCC), .I2C0_SDA_F2H_SCP(VCC), .I2C1_BCLK(VCC)
        , .I2C1_SCL_F2H_SCP(VCC), .I2C1_SDA_F2H_SCP(VCC), .MDIF(VCC), 
        .MGPIO0A_F2H_GPIN(VCC), .MGPIO10A_F2H_GPIN(VCC), 
        .MGPIO11A_F2H_GPIN(VCC), .MGPIO11B_F2H_GPIN(VCC), 
        .MGPIO12A_F2H_GPIN(VCC), .MGPIO13A_F2H_GPIN(VCC), 
        .MGPIO14A_F2H_GPIN(VCC), .MGPIO15A_F2H_GPIN(VCC), 
        .MGPIO16A_F2H_GPIN(VCC), .MGPIO17B_F2H_GPIN(VCC), 
        .MGPIO18B_F2H_GPIN(VCC), .MGPIO19B_F2H_GPIN(VCC), 
        .MGPIO1A_F2H_GPIN(VCC), .MGPIO20B_F2H_GPIN(VCC), 
        .MGPIO21B_F2H_GPIN(VCC), .MGPIO22B_F2H_GPIN(VCC), 
        .MGPIO24B_F2H_GPIN(VCC), .MGPIO25B_F2H_GPIN(VCC), 
        .MGPIO26B_F2H_GPIN(VCC), .MGPIO27B_F2H_GPIN(VCC), 
        .MGPIO28B_F2H_GPIN(VCC), .MGPIO29B_F2H_GPIN(VCC), 
        .MGPIO2A_F2H_GPIN(VCC), .MGPIO30B_F2H_GPIN(VCC), 
        .MGPIO31B_F2H_GPIN(VCC), .MGPIO3A_F2H_GPIN(VCC), 
        .MGPIO4A_F2H_GPIN(VCC), .MGPIO5A_F2H_GPIN(VCC), 
        .MGPIO6A_F2H_GPIN(VCC), .MGPIO7A_F2H_GPIN(VCC), 
        .MGPIO8A_F2H_GPIN(VCC), .MGPIO9A_F2H_GPIN(VCC), 
        .MMUART0_CTS_F2H_SCP(VCC), .MMUART0_DCD_F2H_SCP(VCC), 
        .MMUART0_DSR_F2H_SCP(VCC), .MMUART0_DTR_F2H_SCP(VCC), 
        .MMUART0_RI_F2H_SCP(VCC), .MMUART0_RTS_F2H_SCP(VCC), 
        .MMUART0_RXD_F2H_SCP(VCC), .MMUART0_SCK_F2H_SCP(VCC), 
        .MMUART0_TXD_F2H_SCP(VCC), .MMUART1_CTS_F2H_SCP(VCC), 
        .MMUART1_DCD_F2H_SCP(VCC), .MMUART1_DSR_F2H_SCP(VCC), 
        .MMUART1_RI_F2H_SCP(VCC), .MMUART1_RTS_F2H_SCP(VCC), 
        .MMUART1_RXD_F2H_SCP(VCC), .MMUART1_SCK_F2H_SCP(VCC), 
        .MMUART1_TXD_F2H_SCP(VCC), .PER2_FABRIC_PRDATA({VCC, VCC, VCC, 
        VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, 
        VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, 
        VCC, VCC, VCC, VCC, VCC}), .PER2_FABRIC_PREADY(VCC), 
        .PER2_FABRIC_PSLVERR(VCC), .RCGF({VCC, VCC, VCC, VCC, VCC, VCC, 
        VCC, VCC, VCC, VCC}), .RX_CLKPF(MAC_MII_RX_CLK), .RX_DVF(
        MAC_MII_RX_DV), .RX_ERRF(MAC_MII_RX_ER), .RX_EV(VCC), .RXDF({
        VCC, VCC, VCC, VCC, MAC_MII_RXD[3], MAC_MII_RXD[2], 
        MAC_MII_RXD[1], MAC_MII_RXD[0]}), .SLEEPHOLDREQ(GND), 
        .SMBALERT_NI0(VCC), .SMBALERT_NI1(VCC), .SMBSUS_NI0(VCC), 
        .SMBSUS_NI1(VCC), .SPI0_CLK_IN(VCC), .SPI0_SDI_F2H_SCP(VCC), 
        .SPI0_SDO_F2H_SCP(VCC), .SPI0_SS0_F2H_SCP(VCC), 
        .SPI0_SS1_F2H_SCP(VCC), .SPI0_SS2_F2H_SCP(VCC), 
        .SPI0_SS3_F2H_SCP(VCC), .SPI1_CLK_IN(VCC), .SPI1_SDI_F2H_SCP(
        VCC), .SPI1_SDO_F2H_SCP(VCC), .SPI1_SS0_F2H_SCP(VCC), 
        .SPI1_SS1_F2H_SCP(VCC), .SPI1_SS2_F2H_SCP(VCC), 
        .SPI1_SS3_F2H_SCP(VCC), .TX_CLKPF(MAC_MII_TX_CLK), 
        .USER_MSS_GPIO_RESET_N(VCC), .USER_MSS_RESET_N(VCC), .XCLK_FAB(
        VCC), .CLK_BASE(MCCC_CLK_BASE), .CLK_MDDR_APB(VCC), 
        .F_ARADDR_HADDR1({VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, 
        VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, 
        VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC}), 
        .F_ARBURST_HTRANS1({GND, GND}), .F_ARID_HSEL1({GND, GND, GND, 
        GND}), .F_ARLEN_HBURST1({GND, GND, GND, GND}), 
        .F_ARLOCK_HMASTLOCK1({GND, GND}), .F_ARSIZE_HSIZE1({GND, GND}), 
        .F_ARVALID_HWRITE1(GND), .F_AWADDR_HADDR0({VCC, VCC, VCC, VCC, 
        VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, 
        VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, 
        VCC, VCC, VCC, VCC}), .F_AWBURST_HTRANS0({GND, GND}), 
        .F_AWID_HSEL0({GND, GND, GND, GND}), .F_AWLEN_HBURST0({GND, 
        GND, GND, GND}), .F_AWLOCK_HMASTLOCK0({GND, GND}), 
        .F_AWSIZE_HSIZE0({GND, GND}), .F_AWVALID_HWRITE0(GND), 
        .F_BREADY(GND), .F_RMW_AXI(GND), .F_RREADY(GND), 
        .F_WDATA_HWDATA01({VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, 
        VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, 
        VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, 
        VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, 
        VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, 
        VCC, VCC, VCC, VCC, VCC, VCC, VCC}), .F_WID_HREADY01({GND, GND, 
        GND, GND}), .F_WLAST(GND), .F_WSTRB({GND, GND, GND, GND, GND, 
        GND, GND, GND}), .F_WVALID(GND), .FPGA_MDDR_ARESET_N(VCC), 
        .MDDR_FABRIC_PADDR({VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, 
        VCC}), .MDDR_FABRIC_PENABLE(VCC), .MDDR_FABRIC_PSEL(VCC), 
        .MDDR_FABRIC_PWDATA({VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC, 
        VCC, VCC, VCC, VCC, VCC, VCC, VCC, VCC}), .MDDR_FABRIC_PWRITE(
        VCC), .PRESET_N(GND), .CAN_RXBUS_USBA_DATA1_MGPIO3A_IN(GND), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN(GND), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_IN(GND), .DM_IN({GND, 
        MDDR_DM_RDQS_1_PAD_Y, MDDR_DM_RDQS_0_PAD_Y}), .DRAM_DQ_IN({GND, 
        GND, MDDR_DQ_15_PAD_Y, MDDR_DQ_14_PAD_Y, MDDR_DQ_13_PAD_Y, 
        MDDR_DQ_12_PAD_Y, MDDR_DQ_11_PAD_Y, MDDR_DQ_10_PAD_Y, 
        MDDR_DQ_9_PAD_Y, MDDR_DQ_8_PAD_Y, MDDR_DQ_7_PAD_Y, 
        MDDR_DQ_6_PAD_Y, MDDR_DQ_5_PAD_Y, MDDR_DQ_4_PAD_Y, 
        MDDR_DQ_3_PAD_Y, MDDR_DQ_2_PAD_Y, MDDR_DQ_1_PAD_Y, 
        MDDR_DQ_0_PAD_Y}), .DRAM_DQS_IN({GND, MDDR_DQS_1_PAD_Y, 
        MDDR_DQS_0_PAD_Y}), .DRAM_FIFO_WE_IN({GND, 
        MDDR_DQS_TMATCH_0_IN_PAD_Y}), .I2C0_SCL_USBC_DATA1_MGPIO31B_IN(
        I2C_0_SCL_PAD_Y), .I2C0_SDA_USBC_DATA0_MGPIO30B_IN(
        I2C_0_SDA_PAD_Y), .I2C1_SCL_USBA_DATA4_MGPIO1A_IN(
        I2C_1_SCL_PAD_Y), .I2C1_SDA_USBA_DATA3_MGPIO0A_IN(
        I2C_1_SDA_PAD_Y), .MMUART0_CTS_USBC_DATA7_MGPIO19B_IN(GND), 
        .MMUART0_DCD_MGPIO22B_IN(GND), .MMUART0_DSR_MGPIO20B_IN(GND), 
        .MMUART0_DTR_USBC_DATA6_MGPIO18B_IN(GND), 
        .MMUART0_RI_MGPIO21B_IN(GND), 
        .MMUART0_RTS_USBC_DATA5_MGPIO17B_IN(GND), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_IN(MMUART_0_RXD_PAD_Y), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_IN(GND), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_IN(GND), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_IN(MMUART_1_RXD_PAD_Y), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_IN(GND), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_IN(GND), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN(USB_ULPI_XCLK_PAD_Y), 
        .RGMII_MDC_RMII_MDC_IN(GND), 
        .RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN(USB_ULPI_DATA_7_PAD_Y), 
        .RGMII_RX_CLK_IN(GND), .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN(
        USB_ULPI_DATA_2_PAD_Y), .RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN(
        USB_ULPI_DATA_0_PAD_Y), .RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN(
        USB_ULPI_DATA_1_PAD_Y), .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN(
        USB_ULPI_DATA_3_PAD_Y), .RGMII_RXD3_USBB_DATA4_IN(
        USB_ULPI_DATA_4_PAD_Y), .RGMII_TX_CLK_IN(GND), 
        .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN(USB_ULPI_NXT_PAD_Y), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_IN(USB_ULPI_DIR_PAD_Y), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_IN(GND), 
        .RGMII_TXD2_USBB_DATA5_IN(USB_ULPI_DATA_5_PAD_Y), 
        .RGMII_TXD3_USBB_DATA6_IN(USB_ULPI_DATA_6_PAD_Y), 
        .SPI0_SCK_USBA_XCLK_IN(SPI_0_CLK_PAD_Y), 
        .SPI0_SDI_USBA_DIR_MGPIO5A_IN(SPI_0_DI_PAD_Y), 
        .SPI0_SDO_USBA_STP_MGPIO6A_IN(GND), 
        .SPI0_SS0_USBA_NXT_MGPIO7A_IN(SPI_0_SS0_PAD_Y), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_IN(GND), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_IN(GND), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_IN(GND), .SPI1_SCK_IN(
        SPI_1_CLK_PAD_Y), .SPI1_SDI_MGPIO11A_IN(SPI_1_DI_PAD_Y), 
        .SPI1_SDO_MGPIO12A_IN(GND), .SPI1_SS0_MGPIO13A_IN(
        SPI_1_SS0_PAD_Y), .SPI1_SS1_MGPIO14A_IN(GND), 
        .SPI1_SS2_MGPIO15A_IN(GND), .SPI1_SS3_MGPIO16A_IN(GND), 
        .SPI1_SS4_MGPIO17A_IN(GND), .SPI1_SS5_MGPIO18A_IN(GND), 
        .SPI1_SS6_MGPIO23A_IN(GND), .SPI1_SS7_MGPIO24A_IN(GND), 
        .USBC_XCLK_IN(GND), .CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT(
        CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT(
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT(
        CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT), .DRAM_ADDR({
        DRAM_ADDR_net_0[15], DRAM_ADDR_net_0[14], DRAM_ADDR_net_0[13], 
        DRAM_ADDR_net_0[12], DRAM_ADDR_net_0[11], DRAM_ADDR_net_0[10], 
        DRAM_ADDR_net_0[9], DRAM_ADDR_net_0[8], DRAM_ADDR_net_0[7], 
        DRAM_ADDR_net_0[6], DRAM_ADDR_net_0[5], DRAM_ADDR_net_0[4], 
        DRAM_ADDR_net_0[3], DRAM_ADDR_net_0[2], DRAM_ADDR_net_0[1], 
        DRAM_ADDR_net_0[0]}), .DRAM_BA({DRAM_BA_net_0[2], 
        DRAM_BA_net_0[1], DRAM_BA_net_0[0]}), .DRAM_CASN(
        MSS_ADLIB_INST_DRAM_CASN), .DRAM_CKE(MSS_ADLIB_INST_DRAM_CKE), 
        .DRAM_CLK(MSS_ADLIB_INST_DRAM_CLK), .DRAM_CSN(
        MSS_ADLIB_INST_DRAM_CSN), .DRAM_DM_RDQS_OUT({
        DRAM_DM_RDQS_OUT_net_0[2], DRAM_DM_RDQS_OUT_net_0[1], 
        DRAM_DM_RDQS_OUT_net_0[0]}), .DRAM_DQ_OUT({
        DRAM_DQ_OUT_net_0[17], DRAM_DQ_OUT_net_0[16], 
        DRAM_DQ_OUT_net_0[15], DRAM_DQ_OUT_net_0[14], 
        DRAM_DQ_OUT_net_0[13], DRAM_DQ_OUT_net_0[12], 
        DRAM_DQ_OUT_net_0[11], DRAM_DQ_OUT_net_0[10], 
        DRAM_DQ_OUT_net_0[9], DRAM_DQ_OUT_net_0[8], 
        DRAM_DQ_OUT_net_0[7], DRAM_DQ_OUT_net_0[6], 
        DRAM_DQ_OUT_net_0[5], DRAM_DQ_OUT_net_0[4], 
        DRAM_DQ_OUT_net_0[3], DRAM_DQ_OUT_net_0[2], 
        DRAM_DQ_OUT_net_0[1], DRAM_DQ_OUT_net_0[0]}), .DRAM_DQS_OUT({
        DRAM_DQS_OUT_net_0[2], DRAM_DQS_OUT_net_0[1], 
        DRAM_DQS_OUT_net_0[0]}), .DRAM_FIFO_WE_OUT({
        DRAM_FIFO_WE_OUT_net_0[1], DRAM_FIFO_WE_OUT_net_0[0]}), 
        .DRAM_ODT(MSS_ADLIB_INST_DRAM_ODT), .DRAM_RASN(
        MSS_ADLIB_INST_DRAM_RASN), .DRAM_RSTN(MSS_ADLIB_INST_DRAM_RSTN)
        , .DRAM_WEN(MSS_ADLIB_INST_DRAM_WEN), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_OUT(
        MSS_ADLIB_INST_I2C0_SCL_USBC_DATA1_MGPIO31B_OUT), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_OUT(
        MSS_ADLIB_INST_I2C0_SDA_USBC_DATA0_MGPIO30B_OUT), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_OUT(
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OUT), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_OUT(
        MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OUT), 
        .MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT(
        MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT), 
        .MMUART0_DCD_MGPIO22B_OUT(MMUART0_DCD_MGPIO22B_OUT), 
        .MMUART0_DSR_MGPIO20B_OUT(MMUART0_DSR_MGPIO20B_OUT), 
        .MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT(
        MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT), .MMUART0_RI_MGPIO21B_OUT(
        MMUART0_RI_MGPIO21B_OUT), .MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT(
        MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_OUT(
        MMUART0_RXD_USBC_STP_MGPIO28B_OUT), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_OUT(
        MMUART0_SCK_USBC_NXT_MGPIO29B_OUT), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_OUT(
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OUT), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT(
        MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT(
        MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT(
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT(
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT), .RGMII_MDC_RMII_MDC_OUT(
        RGMII_MDC_RMII_MDC_OUT), .RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT(
        MSS_ADLIB_INST_RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT), 
        .RGMII_RX_CLK_OUT(RGMII_RX_CLK_OUT), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT(
        MSS_ADLIB_INST_RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT(
        MSS_ADLIB_INST_RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT(
        MSS_ADLIB_INST_RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT(
        MSS_ADLIB_INST_RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT), 
        .RGMII_RXD3_USBB_DATA4_OUT(
        MSS_ADLIB_INST_RGMII_RXD3_USBB_DATA4_OUT), .RGMII_TX_CLK_OUT(
        RGMII_TX_CLK_OUT), .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT(
        RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT(
        RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_OUT(
        MSS_ADLIB_INST_RGMII_TXD1_RMII_TXD1_USBB_STP_OUT), 
        .RGMII_TXD2_USBB_DATA5_OUT(
        MSS_ADLIB_INST_RGMII_TXD2_USBB_DATA5_OUT), 
        .RGMII_TXD3_USBB_DATA6_OUT(
        MSS_ADLIB_INST_RGMII_TXD3_USBB_DATA6_OUT), 
        .SPI0_SCK_USBA_XCLK_OUT(MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OUT), 
        .SPI0_SDI_USBA_DIR_MGPIO5A_OUT(SPI0_SDI_USBA_DIR_MGPIO5A_OUT), 
        .SPI0_SDO_USBA_STP_MGPIO6A_OUT(
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OUT), 
        .SPI0_SS0_USBA_NXT_MGPIO7A_OUT(
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OUT), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_OUT(
        SPI0_SS1_USBA_DATA5_MGPIO8A_OUT), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_OUT(
        SPI0_SS2_USBA_DATA6_MGPIO9A_OUT), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_OUT(
        SPI0_SS3_USBA_DATA7_MGPIO10A_OUT), .SPI1_SCK_OUT(
        MSS_ADLIB_INST_SPI1_SCK_OUT), .SPI1_SDI_MGPIO11A_OUT(
        SPI1_SDI_MGPIO11A_OUT), .SPI1_SDO_MGPIO12A_OUT(
        MSS_ADLIB_INST_SPI1_SDO_MGPIO12A_OUT), .SPI1_SS0_MGPIO13A_OUT(
        MSS_ADLIB_INST_SPI1_SS0_MGPIO13A_OUT), .SPI1_SS1_MGPIO14A_OUT(
        SPI1_SS1_MGPIO14A_OUT), .SPI1_SS2_MGPIO15A_OUT(
        SPI1_SS2_MGPIO15A_OUT), .SPI1_SS3_MGPIO16A_OUT(
        SPI1_SS3_MGPIO16A_OUT), .SPI1_SS4_MGPIO17A_OUT(
        SPI1_SS4_MGPIO17A_OUT), .SPI1_SS5_MGPIO18A_OUT(
        SPI1_SS5_MGPIO18A_OUT), .SPI1_SS6_MGPIO23A_OUT(
        SPI1_SS6_MGPIO23A_OUT), .SPI1_SS7_MGPIO24A_OUT(
        SPI1_SS7_MGPIO24A_OUT), .USBC_XCLK_OUT(USBC_XCLK_OUT), 
        .CAN_RXBUS_USBA_DATA1_MGPIO3A_OE(
        CAN_RXBUS_USBA_DATA1_MGPIO3A_OE), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE(
        CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_OE(
        CAN_TXBUS_USBA_DATA0_MGPIO2A_OE), .DM_OE({DM_OE_net_0[2], 
        DM_OE_net_0[1], DM_OE_net_0[0]}), .DRAM_DQ_OE({
        DRAM_DQ_OE_net_0[17], DRAM_DQ_OE_net_0[16], 
        DRAM_DQ_OE_net_0[15], DRAM_DQ_OE_net_0[14], 
        DRAM_DQ_OE_net_0[13], DRAM_DQ_OE_net_0[12], 
        DRAM_DQ_OE_net_0[11], DRAM_DQ_OE_net_0[10], 
        DRAM_DQ_OE_net_0[9], DRAM_DQ_OE_net_0[8], DRAM_DQ_OE_net_0[7], 
        DRAM_DQ_OE_net_0[6], DRAM_DQ_OE_net_0[5], DRAM_DQ_OE_net_0[4], 
        DRAM_DQ_OE_net_0[3], DRAM_DQ_OE_net_0[2], DRAM_DQ_OE_net_0[1], 
        DRAM_DQ_OE_net_0[0]}), .DRAM_DQS_OE({DRAM_DQS_OE_net_0[2], 
        DRAM_DQS_OE_net_0[1], DRAM_DQS_OE_net_0[0]}), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_OE(
        MSS_ADLIB_INST_I2C0_SCL_USBC_DATA1_MGPIO31B_OE), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_OE(
        MSS_ADLIB_INST_I2C0_SDA_USBC_DATA0_MGPIO30B_OE), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_OE(
        MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OE), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_OE(
        MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OE), 
        .MMUART0_CTS_USBC_DATA7_MGPIO19B_OE(
        MMUART0_CTS_USBC_DATA7_MGPIO19B_OE), .MMUART0_DCD_MGPIO22B_OE(
        MMUART0_DCD_MGPIO22B_OE), .MMUART0_DSR_MGPIO20B_OE(
        MMUART0_DSR_MGPIO20B_OE), .MMUART0_DTR_USBC_DATA6_MGPIO18B_OE(
        MMUART0_DTR_USBC_DATA6_MGPIO18B_OE), .MMUART0_RI_MGPIO21B_OE(
        MMUART0_RI_MGPIO21B_OE), .MMUART0_RTS_USBC_DATA5_MGPIO17B_OE(
        MMUART0_RTS_USBC_DATA5_MGPIO17B_OE), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_OE(
        MMUART0_RXD_USBC_STP_MGPIO28B_OE), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_OE(
        MMUART0_SCK_USBC_NXT_MGPIO29B_OE), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_OE(
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OE), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_OE(
        MMUART1_RXD_USBC_DATA3_MGPIO26B_OE), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_OE(
        MMUART1_SCK_USBC_DATA4_MGPIO25B_OE), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_OE(
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OE), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE(
        RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE), .RGMII_MDC_RMII_MDC_OE(
        RGMII_MDC_RMII_MDC_OE), .RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE(
        MSS_ADLIB_INST_RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE), 
        .RGMII_RX_CLK_OE(RGMII_RX_CLK_OE), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE(
        MSS_ADLIB_INST_RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE(
        MSS_ADLIB_INST_RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE(
        MSS_ADLIB_INST_RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE(
        MSS_ADLIB_INST_RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE), 
        .RGMII_RXD3_USBB_DATA4_OE(
        MSS_ADLIB_INST_RGMII_RXD3_USBB_DATA4_OE), .RGMII_TX_CLK_OE(
        RGMII_TX_CLK_OE), .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE(
        RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_OE(
        RGMII_TXD0_RMII_TXD0_USBB_DIR_OE), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_OE(
        MSS_ADLIB_INST_RGMII_TXD1_RMII_TXD1_USBB_STP_OE), 
        .RGMII_TXD2_USBB_DATA5_OE(
        MSS_ADLIB_INST_RGMII_TXD2_USBB_DATA5_OE), 
        .RGMII_TXD3_USBB_DATA6_OE(
        MSS_ADLIB_INST_RGMII_TXD3_USBB_DATA6_OE), 
        .SPI0_SCK_USBA_XCLK_OE(MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OE), 
        .SPI0_SDI_USBA_DIR_MGPIO5A_OE(SPI0_SDI_USBA_DIR_MGPIO5A_OE), 
        .SPI0_SDO_USBA_STP_MGPIO6A_OE(
        MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OE), 
        .SPI0_SS0_USBA_NXT_MGPIO7A_OE(
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OE), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_OE(SPI0_SS1_USBA_DATA5_MGPIO8A_OE)
        , .SPI0_SS2_USBA_DATA6_MGPIO9A_OE(
        SPI0_SS2_USBA_DATA6_MGPIO9A_OE), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_OE(
        SPI0_SS3_USBA_DATA7_MGPIO10A_OE), .SPI1_SCK_OE(
        MSS_ADLIB_INST_SPI1_SCK_OE), .SPI1_SDI_MGPIO11A_OE(
        SPI1_SDI_MGPIO11A_OE), .SPI1_SDO_MGPIO12A_OE(
        MSS_ADLIB_INST_SPI1_SDO_MGPIO12A_OE), .SPI1_SS0_MGPIO13A_OE(
        MSS_ADLIB_INST_SPI1_SS0_MGPIO13A_OE), .SPI1_SS1_MGPIO14A_OE(
        SPI1_SS1_MGPIO14A_OE), .SPI1_SS2_MGPIO15A_OE(
        SPI1_SS2_MGPIO15A_OE), .SPI1_SS3_MGPIO16A_OE(
        SPI1_SS3_MGPIO16A_OE), .SPI1_SS4_MGPIO17A_OE(
        SPI1_SS4_MGPIO17A_OE), .SPI1_SS5_MGPIO18A_OE(
        SPI1_SS5_MGPIO18A_OE), .SPI1_SS6_MGPIO23A_OE(
        SPI1_SS6_MGPIO23A_OE), .SPI1_SS7_MGPIO24A_OE(
        SPI1_SS7_MGPIO24A_OE), .USBC_XCLK_OE(USBC_XCLK_OE));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_RAS_N_PAD (.D(
        MSS_ADLIB_INST_DRAM_RASN), .PAD(MDDR_RAS_N));
    BIBUF #( .IOSTD("") )  SPI_0_CLK_PAD (.PAD(SPI_0_CLK), .D(
        MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OUT), .E(
        MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OE), .Y(SPI_0_CLK_PAD_Y));
    BIBUF #( .IOSTD("") )  USB_ULPI_DATA_1_PAD (.PAD(USB_ULPI_DATA[1]), 
        .D(MSS_ADLIB_INST_RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT), .E(
        MSS_ADLIB_INST_RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE), .Y(
        USB_ULPI_DATA_1_PAD_Y));
    BIBUF #( .IOSTD("SSTL18I") )  MDDR_DQ_4_PAD (.PAD(MDDR_DQ[4]), .D(
        DRAM_DQ_OUT_net_0[4]), .E(DRAM_DQ_OE_net_0[4]), .Y(
        MDDR_DQ_4_PAD_Y));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_ADDR_10_PAD (.D(
        DRAM_ADDR_net_0[10]), .PAD(MDDR_ADDR[10]));
    BIBUF #( .IOSTD("") )  I2C_0_SDA_PAD (.PAD(I2C_0_SDA), .D(
        MSS_ADLIB_INST_I2C0_SDA_USBC_DATA0_MGPIO30B_OUT), .E(
        MSS_ADLIB_INST_I2C0_SDA_USBC_DATA0_MGPIO30B_OE), .Y(
        I2C_0_SDA_PAD_Y));
    INBUF #( .IOSTD("SSTL18I") )  MDDR_DQS_TMATCH_0_IN_PAD (.PAD(
        MDDR_DQS_TMATCH_0_IN), .Y(MDDR_DQS_TMATCH_0_IN_PAD_Y));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_CS_N_PAD (.D(
        MSS_ADLIB_INST_DRAM_CSN), .PAD(MDDR_CS_N));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_ADDR_4_PAD (.D(
        DRAM_ADDR_net_0[4]), .PAD(MDDR_ADDR[4]));
    GND GND_Z (.Y(GND));
    VCC VCC_Z (.Y(VCC));
    BIBUF #( .IOSTD("") )  USB_ULPI_DATA_5_PAD (.PAD(USB_ULPI_DATA[5]), 
        .D(MSS_ADLIB_INST_RGMII_TXD2_USBB_DATA5_OUT), .E(
        MSS_ADLIB_INST_RGMII_TXD2_USBB_DATA5_OE), .Y(
        USB_ULPI_DATA_5_PAD_Y));
    BIBUF #( .IOSTD("") )  SPI_0_SS0_PAD (.PAD(SPI_0_SS0), .D(
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OUT), .E(
        MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OE), .Y(
        SPI_0_SS0_PAD_Y));
    BIBUF #( .IOSTD("SSTL18I") )  MDDR_DQ_7_PAD (.PAD(MDDR_DQ[7]), .D(
        DRAM_DQ_OUT_net_0[7]), .E(DRAM_DQ_OE_net_0[7]), .Y(
        MDDR_DQ_7_PAD_Y));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_WE_N_PAD (.D(
        MSS_ADLIB_INST_DRAM_WEN), .PAD(MDDR_WE_N));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_ADDR_8_PAD (.D(
        DRAM_ADDR_net_0[8]), .PAD(MDDR_ADDR[8]));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_ADDR_15_PAD (.D(
        DRAM_ADDR_net_0[15]), .PAD(MDDR_ADDR[15]));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_ADDR_0_PAD (.D(
        DRAM_ADDR_net_0[0]), .PAD(MDDR_ADDR[0]));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_ADDR_1_PAD (.D(
        DRAM_ADDR_net_0[1]), .PAD(MDDR_ADDR[1]));
    BIBUF #( .IOSTD("SSTL18I") )  MDDR_DQ_13_PAD (.PAD(MDDR_DQ[13]), 
        .D(DRAM_DQ_OUT_net_0[13]), .E(DRAM_DQ_OE_net_0[13]), .Y(
        MDDR_DQ_13_PAD_Y));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_ADDR_3_PAD (.D(
        DRAM_ADDR_net_0[3]), .PAD(MDDR_ADDR[3]));
    INBUF #( .IOSTD("") )  MMUART_1_RXD_PAD (.PAD(MMUART_1_RXD), .Y(
        MMUART_1_RXD_PAD_Y));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_BA_0_PAD (.D(DRAM_BA_net_0[0]), 
        .PAD(MDDR_BA[0]));
    BIBUF #( .IOSTD("SSTL18I") )  MDDR_DQ_6_PAD (.PAD(MDDR_DQ[6]), .D(
        DRAM_DQ_OUT_net_0[6]), .E(DRAM_DQ_OE_net_0[6]), .Y(
        MDDR_DQ_6_PAD_Y));
    OUTBUF_DIFF #( .IOSTD("SSTL18I") )  MDDR_CLK_PAD (.D(
        MSS_ADLIB_INST_DRAM_CLK), .PADP(MDDR_CLK), .PADN(MDDR_CLK_N));
    BIBUF #( .IOSTD("SSTL18I") )  MDDR_DQ_14_PAD (.PAD(MDDR_DQ[14]), 
        .D(DRAM_DQ_OUT_net_0[14]), .E(DRAM_DQ_OE_net_0[14]), .Y(
        MDDR_DQ_14_PAD_Y));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_DQS_TMATCH_0_OUT_PAD (.D(
        DRAM_FIFO_WE_OUT_net_0[0]), .PAD(MDDR_DQS_TMATCH_0_OUT));
    INBUF #( .IOSTD("") )  USB_ULPI_NXT_PAD (.PAD(USB_ULPI_NXT), .Y(
        USB_ULPI_NXT_PAD_Y));
    OUTBUF #( .IOSTD("SSTL18I") )  MDDR_BA_1_PAD (.D(DRAM_BA_net_0[1]), 
        .PAD(MDDR_BA[1]));
    BIBUF #( .IOSTD("") )  USB_ULPI_DATA_6_PAD (.PAD(USB_ULPI_DATA[6]), 
        .D(MSS_ADLIB_INST_RGMII_TXD3_USBB_DATA6_OUT), .E(
        MSS_ADLIB_INST_RGMII_TXD3_USBB_DATA6_OE), .Y(
        USB_ULPI_DATA_6_PAD_Y));
    BIBUF #( .IOSTD("") )  SPI_1_CLK_PAD (.PAD(SPI_1_CLK), .D(
        MSS_ADLIB_INST_SPI1_SCK_OUT), .E(MSS_ADLIB_INST_SPI1_SCK_OE), 
        .Y(SPI_1_CLK_PAD_Y));
    BIBUF #( .IOSTD("SSTL18I") )  MDDR_DQ_5_PAD (.PAD(MDDR_DQ[5]), .D(
        DRAM_DQ_OUT_net_0[5]), .E(DRAM_DQ_OE_net_0[5]), .Y(
        MDDR_DQ_5_PAD_Y));
    
endmodule


module SF2Project(
       MAC_MII_COL,
       MAC_MII_CRS,
       MAC_MII_RXD,
       MAC_MII_RX_CLK,
       MAC_MII_RX_DV,
       MAC_MII_RX_ER,
       MAC_MII_TX_CLK,
       MCCC_CLK_BASE,
       MDDR_DQS_TMATCH_0_IN,
       MMUART_0_RXD,
       MMUART_1_RXD,
       SPI_0_DI,
       SPI_1_DI,
       USB_ULPI_DIR,
       USB_ULPI_NXT,
       USB_ULPI_XCLK,
       MAC_MII_TXD,
       MAC_MII_TX_EN,
       MAC_MII_TX_ER,
       MDDR_ADDR,
       MDDR_BA,
       MDDR_CAS_N,
       MDDR_CKE,
       MDDR_CLK,
       MDDR_CLK_N,
       MDDR_CS_N,
       MDDR_DQS_TMATCH_0_OUT,
       MDDR_ODT,
       MDDR_RAS_N,
       MDDR_RESET_N,
       MDDR_WE_N,
       MMUART_0_TXD,
       MMUART_1_TXD,
       SPI_0_DO,
       SPI_1_DO,
       USB_ULPI_STP,
       I2C_0_SCL,
       I2C_0_SDA,
       I2C_1_SCL,
       I2C_1_SDA,
       MDDR_DM_RDQS,
       MDDR_DQ,
       MDDR_DQS,
       MDDR_DQS_N,
       SPI_0_CLK,
       SPI_0_SS0,
       SPI_1_CLK,
       SPI_1_SS0,
       USB_ULPI_DATA
    );
input  MAC_MII_COL;
input  MAC_MII_CRS;
input  [3:0] MAC_MII_RXD;
input  MAC_MII_RX_CLK;
input  MAC_MII_RX_DV;
input  MAC_MII_RX_ER;
input  MAC_MII_TX_CLK;
input  MCCC_CLK_BASE;
input  MDDR_DQS_TMATCH_0_IN;
input  MMUART_0_RXD;
input  MMUART_1_RXD;
input  SPI_0_DI;
input  SPI_1_DI;
input  USB_ULPI_DIR;
input  USB_ULPI_NXT;
input  USB_ULPI_XCLK;
output [3:0] MAC_MII_TXD;
output MAC_MII_TX_EN;
output MAC_MII_TX_ER;
output [15:0] MDDR_ADDR;
output [2:0] MDDR_BA;
output MDDR_CAS_N;
output MDDR_CKE;
output MDDR_CLK;
output MDDR_CLK_N;
output MDDR_CS_N;
output MDDR_DQS_TMATCH_0_OUT;
output MDDR_ODT;
output MDDR_RAS_N;
output MDDR_RESET_N;
output MDDR_WE_N;
output MMUART_0_TXD;
output MMUART_1_TXD;
output SPI_0_DO;
output SPI_1_DO;
output USB_ULPI_STP;
inout  I2C_0_SCL;
inout  I2C_0_SDA;
inout  I2C_1_SCL;
inout  I2C_1_SDA;
inout  [1:0] MDDR_DM_RDQS;
inout  [15:0] MDDR_DQ;
inout  [1:0] MDDR_DQS;
inout  [1:0] MDDR_DQS_N;
inout  SPI_0_CLK;
inout  SPI_0_SS0;
inout  SPI_1_CLK;
inout  SPI_1_SS0;
inout  [7:0] USB_ULPI_DATA;

    wire GND, VCC;
    
    SF2Project_MSS SF2Project_MSS_0 (.MDDR_DQS({MDDR_DQS[1], 
        MDDR_DQS[0]}), .MDDR_DQS_N({MDDR_DQS_N[1], MDDR_DQS_N[0]}), 
        .MAC_MII_RXD({MAC_MII_RXD[3], MAC_MII_RXD[2], MAC_MII_RXD[1], 
        MAC_MII_RXD[0]}), .MAC_MII_TXD({MAC_MII_TXD[3], MAC_MII_TXD[2], 
        MAC_MII_TXD[1], MAC_MII_TXD[0]}), .MDDR_ADDR({MDDR_ADDR[15], 
        MDDR_ADDR[14], MDDR_ADDR[13], MDDR_ADDR[12], MDDR_ADDR[11], 
        MDDR_ADDR[10], MDDR_ADDR[9], MDDR_ADDR[8], MDDR_ADDR[7], 
        MDDR_ADDR[6], MDDR_ADDR[5], MDDR_ADDR[4], MDDR_ADDR[3], 
        MDDR_ADDR[2], MDDR_ADDR[1], MDDR_ADDR[0]}), .MDDR_BA({
        MDDR_BA[2], MDDR_BA[1], MDDR_BA[0]}), .MDDR_DM_RDQS({
        MDDR_DM_RDQS[1], MDDR_DM_RDQS[0]}), .MDDR_DQ({MDDR_DQ[15], 
        MDDR_DQ[14], MDDR_DQ[13], MDDR_DQ[12], MDDR_DQ[11], 
        MDDR_DQ[10], MDDR_DQ[9], MDDR_DQ[8], MDDR_DQ[7], MDDR_DQ[6], 
        MDDR_DQ[5], MDDR_DQ[4], MDDR_DQ[3], MDDR_DQ[2], MDDR_DQ[1], 
        MDDR_DQ[0]}), .USB_ULPI_DATA({USB_ULPI_DATA[7], 
        USB_ULPI_DATA[6], USB_ULPI_DATA[5], USB_ULPI_DATA[4], 
        USB_ULPI_DATA[3], USB_ULPI_DATA[2], USB_ULPI_DATA[1], 
        USB_ULPI_DATA[0]}), .MDDR_CLK(MDDR_CLK), .MDDR_CLK_N(
        MDDR_CLK_N), .MCCC_CLK_BASE(MCCC_CLK_BASE), .MAC_MII_TX_CLK(
        MAC_MII_TX_CLK), .MAC_MII_RX_ER(MAC_MII_RX_ER), .MAC_MII_RX_DV(
        MAC_MII_RX_DV), .MAC_MII_RX_CLK(MAC_MII_RX_CLK), .MAC_MII_CRS(
        MAC_MII_CRS), .MAC_MII_COL(MAC_MII_COL), .MAC_MII_TX_ER(
        MAC_MII_TX_ER), .MAC_MII_TX_EN(MAC_MII_TX_EN), .I2C_0_SCL(
        I2C_0_SCL), .I2C_0_SDA(I2C_0_SDA), .I2C_1_SCL(I2C_1_SCL), 
        .I2C_1_SDA(I2C_1_SDA), .MDDR_CAS_N(MDDR_CAS_N), .MDDR_CKE(
        MDDR_CKE), .MDDR_CS_N(MDDR_CS_N), .MDDR_DQS_TMATCH_0_IN(
        MDDR_DQS_TMATCH_0_IN), .MDDR_DQS_TMATCH_0_OUT(
        MDDR_DQS_TMATCH_0_OUT), .MDDR_ODT(MDDR_ODT), .MDDR_RAS_N(
        MDDR_RAS_N), .MDDR_RESET_N(MDDR_RESET_N), .MDDR_WE_N(MDDR_WE_N)
        , .MMUART_0_RXD(MMUART_0_RXD), .MMUART_0_TXD(MMUART_0_TXD), 
        .MMUART_1_RXD(MMUART_1_RXD), .MMUART_1_TXD(MMUART_1_TXD), 
        .SPI_0_CLK(SPI_0_CLK), .SPI_0_DI(SPI_0_DI), .SPI_0_DO(SPI_0_DO)
        , .SPI_0_SS0(SPI_0_SS0), .SPI_1_CLK(SPI_1_CLK), .SPI_1_DI(
        SPI_1_DI), .SPI_1_DO(SPI_1_DO), .SPI_1_SS0(SPI_1_SS0), 
        .USB_ULPI_DIR(USB_ULPI_DIR), .USB_ULPI_NXT(USB_ULPI_NXT), 
        .USB_ULPI_STP(USB_ULPI_STP), .USB_ULPI_XCLK(USB_ULPI_XCLK));
    VCC VCC_Z (.Y(VCC));
    GND GND_Z (.Y(GND));
    
endmodule
