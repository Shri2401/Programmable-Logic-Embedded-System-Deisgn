`timescale 1 ns/100 ps
// Version: v12.6 12.900.20.24
// File used only for Simulation


module sdf_IOPAD_TRI(
       PAD,
       D,
       E
    );
output PAD;
input  D;
input  E;

    wire NET_OIN_VDD, NET_EIN_VDD;
    
    IOPAD_TRI_VDDI U_VCCI (.OIN_VDD(NET_OIN_VDD), .EIN_VDD(NET_EIN_VDD)
        , .PAD_P(PAD));
    IOPAD_VDD U_VCCA (.OIN_P(D), .EIN_P(E), .IOUT_VDD(), .OIN_VDD(
        NET_OIN_VDD), .EIN_VDD(NET_EIN_VDD), .IOUT_IN());
    
endmodule


module sdf_IOPADN_BI(
       PAD_P,
       OIN_P,
       EIN_P,
       N2POUT_P
    );
inout  PAD_P;
input  OIN_P;
input  EIN_P;
output N2POUT_P;

    wire NET_IOUT_VDD, NET_IOUT_IN, NET_OIN_VDD, NET_EIN_VDD;
    
    IOPADN_BI_VDDI U_VCCI (.OIN_VDD(NET_OIN_VDD), .EIN_VDD(NET_EIN_VDD)
        , .IOUT_VDD(NET_IOUT_VDD), .PAD_P(PAD_P));
    IOPADN_DELAY U_DELAY (.IOUT_IN(NET_IOUT_IN), .N2POUT_P(N2POUT_P));
    IOPADN_VDD U_VCCA (.OIN_P(OIN_P), .EIN_P(EIN_P), .IOUT_VDD(
        NET_IOUT_VDD), .OIN_VDD(NET_OIN_VDD), .EIN_VDD(NET_EIN_VDD), 
        .IOUT_IN(NET_IOUT_IN));
    
endmodule


module sdf_IOPAD_BI(
       PAD,
       D,
       E,
       Y
    );
inout  PAD;
input  D;
input  E;
output Y;

    wire NET_IOUT_VDD, NET_IOUT_IN, NET_OIN_VDD, NET_EIN_VDD;
    
    IOPAD_BI_VDDI U_VCCI (.OIN_VDD(NET_OIN_VDD), .EIN_VDD(NET_EIN_VDD), 
        .IOUT_VDD(NET_IOUT_VDD), .PAD_P(PAD));
    IOPAD_DELAY U_DELAY (.IOUT_IN(NET_IOUT_IN), .IOUT_P(Y));
    IOPAD_VDD U_VCCA (.OIN_P(D), .EIN_P(E), .IOUT_VDD(NET_IOUT_VDD), 
        .OIN_VDD(NET_OIN_VDD), .EIN_VDD(NET_EIN_VDD), .IOUT_IN(
        NET_IOUT_IN));
    
endmodule


module sdf_IOPADN_TRI(
       PAD_P,
       OIN_P,
       EIN_P
    );
output PAD_P;
input  OIN_P;
input  EIN_P;

    wire NET_OIN_VDD, NET_EIN_VDD;
    
    IOPADN_TRI_VDDI U_VCCI (.OIN_VDD(NET_OIN_VDD), .EIN_VDD(
        NET_EIN_VDD), .PAD_P(PAD_P));
    IOPADN_VDD U_VCCA (.OIN_P(OIN_P), .EIN_P(EIN_P), .IOUT_VDD(), 
        .OIN_VDD(NET_OIN_VDD), .EIN_VDD(NET_EIN_VDD), .IOUT_IN());
    
endmodule


module sdf_IOPAD_IN(
       PAD,
       Y
    );
input  PAD;
output Y;

    wire NET_IOUT_VDD, NET_IOUT_IN, ADLIB_GND;
    wire GND_power_net1;
    assign ADLIB_GND = GND_power_net1;
    
    IOPAD_IN_VDDI U_VCCI (.PAD_P(PAD), .IOUT_VDD(NET_IOUT_VDD));
    IOPAD_DELAY U_DELAY (.IOUT_IN(NET_IOUT_IN), .IOUT_P(Y));
    IOPAD_VDD U_VCCA (.OIN_P(ADLIB_GND), .EIN_P(ADLIB_GND), .IOUT_VDD(
        NET_IOUT_VDD), .OIN_VDD(), .EIN_VDD(), .IOUT_IN(NET_IOUT_IN));
    GND GND_power_inst1 (.Y(GND_power_net1));
    
endmodule


module sdf_IOPADP_BI(
       PAD_P,
       N2PIN_P,
       OIN_P,
       EIN_P,
       IOUT_P
    );
inout  PAD_P;
input  N2PIN_P;
input  OIN_P;
input  EIN_P;
output IOUT_P;

    wire NET_IOUT_VDD, NET_IOUT_IN, NET_OIN_VDD, NET_EIN_VDD;
    
    IOPADP_BI_VDDI U_VCCI (.OIN_VDD(NET_OIN_VDD), .EIN_VDD(NET_EIN_VDD)
        , .N2PIN_P(N2PIN_P), .IOUT_VDD(NET_IOUT_VDD), .PAD_P(PAD_P));
    IOPADP_DELAY U_DELAY (.IOUT_IN(NET_IOUT_IN), .IOUT_P(IOUT_P));
    IOPADP_VDD U_VCCA (.OIN_P(OIN_P), .EIN_P(EIN_P), .IOUT_VDD(
        NET_IOUT_VDD), .OIN_VDD(NET_OIN_VDD), .EIN_VDD(NET_EIN_VDD), 
        .IOUT_IN(NET_IOUT_IN));
    
endmodule


module sdf_IOPADP_TRI(
       PAD_P,
       OIN_P,
       EIN_P
    );
output PAD_P;
input  OIN_P;
input  EIN_P;

    wire NET_OIN_VDD, NET_EIN_VDD;
    
    IOPADP_TRI_VDDI U_VCCI (.OIN_VDD(NET_OIN_VDD), .EIN_VDD(
        NET_EIN_VDD), .PAD_P(PAD_P));
    IOPADP_VDD U_VCCA (.OIN_P(OIN_P), .EIN_P(EIN_P), .IOUT_VDD(), 
        .OIN_VDD(NET_OIN_VDD), .EIN_VDD(NET_EIN_VDD), .IOUT_IN());
    
endmodule


module SF2Project(
       MAC_MII_COL,
       MAC_MII_CRS,
       MAC_MII_RXD,
       MAC_MII_RX_CLK,
       MAC_MII_RX_DV,
       MAC_MII_RX_ER,
       MAC_MII_TX_CLK,
       MCCC_CLK_BASE,
       MDDR_DQS_TMATCH_0_IN,
       MMUART_0_RXD,
       MMUART_1_RXD,
       SPI_0_DI,
       SPI_1_DI,
       USB_ULPI_DIR,
       USB_ULPI_NXT,
       USB_ULPI_XCLK,
       MAC_MII_TXD,
       MAC_MII_TX_EN,
       MAC_MII_TX_ER,
       MDDR_ADDR,
       MDDR_BA,
       MDDR_CAS_N,
       MDDR_CKE,
       MDDR_CLK,
       MDDR_CLK_N,
       MDDR_CS_N,
       MDDR_DQS_TMATCH_0_OUT,
       MDDR_ODT,
       MDDR_RAS_N,
       MDDR_RESET_N,
       MDDR_WE_N,
       MMUART_0_TXD,
       MMUART_1_TXD,
       SPI_0_DO,
       SPI_1_DO,
       USB_ULPI_STP,
       I2C_0_SCL,
       I2C_0_SDA,
       I2C_1_SCL,
       I2C_1_SDA,
       MDDR_DM_RDQS,
       MDDR_DQ,
       MDDR_DQS,
       MDDR_DQS_N,
       SPI_0_CLK,
       SPI_0_SS0,
       SPI_1_CLK,
       SPI_1_SS0,
       USB_ULPI_DATA
    );
input  MAC_MII_COL;
input  MAC_MII_CRS;
input  [3:0] MAC_MII_RXD;
input  MAC_MII_RX_CLK;
input  MAC_MII_RX_DV;
input  MAC_MII_RX_ER;
input  MAC_MII_TX_CLK;
input  MCCC_CLK_BASE;
input  MDDR_DQS_TMATCH_0_IN;
input  MMUART_0_RXD;
input  MMUART_1_RXD;
input  SPI_0_DI;
input  SPI_1_DI;
input  USB_ULPI_DIR;
input  USB_ULPI_NXT;
input  USB_ULPI_XCLK;
output [3:0] MAC_MII_TXD;
output MAC_MII_TX_EN;
output MAC_MII_TX_ER;
output [15:0] MDDR_ADDR;
output [2:0] MDDR_BA;
output MDDR_CAS_N;
output MDDR_CKE;
output MDDR_CLK;
output MDDR_CLK_N;
output MDDR_CS_N;
output MDDR_DQS_TMATCH_0_OUT;
output MDDR_ODT;
output MDDR_RAS_N;
output MDDR_RESET_N;
output MDDR_WE_N;
output MMUART_0_TXD;
output MMUART_1_TXD;
output SPI_0_DO;
output SPI_1_DO;
output USB_ULPI_STP;
inout  I2C_0_SCL;
inout  I2C_0_SDA;
inout  I2C_1_SCL;
inout  I2C_1_SDA;
inout  [1:0] MDDR_DM_RDQS;
inout  [15:0] MDDR_DQ;
inout  [1:0] MDDR_DQS;
inout  [1:0] MDDR_DQS_N;
inout  SPI_0_CLK;
inout  SPI_0_SS0;
inout  SPI_1_CLK;
inout  SPI_1_SS0;
inout  [7:0] USB_ULPI_DATA;

    wire \MAC_MII_RXD[3] , \MAC_MII_RXD[2] , \MAC_MII_RXD[1] , 
        \MAC_MII_RXD[0] , \MAC_MII_TXD[3] , \MAC_MII_TXD[2] , 
        \MAC_MII_TXD[1] , \MAC_MII_TXD[0] , MAC_MII_COL_net_1, 
        MAC_MII_CRS_net_1, MAC_MII_RX_CLK_net_1, MAC_MII_RX_DV_net_1, 
        MAC_MII_RX_ER_net_1, MAC_MII_TX_CLK_net_1, MCCC_CLK_BASE_net_1, 
        MAC_MII_TX_EN_net_1, MAC_MII_TX_ER_net_1, 
        \SF2Project_MSS_0/DRAM_FIFO_WE_OUT_net_0[0] , 
        \SF2Project_MSS_0/DRAM_DQ_OUT_net_0[15] , 
        \SF2Project_MSS_0/DRAM_DQ_OUT_net_0[14] , 
        \SF2Project_MSS_0/DRAM_DQ_OUT_net_0[13] , 
        \SF2Project_MSS_0/DRAM_DQ_OUT_net_0[12] , 
        \SF2Project_MSS_0/DRAM_DQ_OUT_net_0[11] , 
        \SF2Project_MSS_0/DRAM_DQ_OUT_net_0[10] , 
        \SF2Project_MSS_0/DRAM_DQ_OUT_net_0[9] , 
        \SF2Project_MSS_0/DRAM_DQ_OUT_net_0[8] , 
        \SF2Project_MSS_0/DRAM_DQ_OUT_net_0[7] , 
        \SF2Project_MSS_0/DRAM_DQ_OUT_net_0[6] , 
        \SF2Project_MSS_0/DRAM_DQ_OUT_net_0[5] , 
        \SF2Project_MSS_0/DRAM_DQ_OUT_net_0[4] , 
        \SF2Project_MSS_0/DRAM_DQ_OUT_net_0[3] , 
        \SF2Project_MSS_0/DRAM_DQ_OUT_net_0[2] , 
        \SF2Project_MSS_0/DRAM_DQ_OUT_net_0[1] , 
        \SF2Project_MSS_0/DRAM_DQ_OUT_net_0[0] , 
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[15] , 
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[14] , 
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[13] , 
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[12] , 
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[11] , 
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[10] , 
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[9] , 
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[8] , 
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[7] , 
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[6] , 
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[5] , 
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[4] , 
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[3] , 
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[2] , 
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[1] , 
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[0] , 
        \SF2Project_MSS_0/DRAM_DM_RDQS_OUT_net_0[1] , 
        \SF2Project_MSS_0/DRAM_DM_RDQS_OUT_net_0[0] , 
        \SF2Project_MSS_0/DM_OE_net_0[1] , 
        \SF2Project_MSS_0/DM_OE_net_0[0] , 
        \SF2Project_MSS_0/DRAM_BA_net_0[2] , 
        \SF2Project_MSS_0/DRAM_BA_net_0[1] , 
        \SF2Project_MSS_0/DRAM_BA_net_0[0] , 
        \SF2Project_MSS_0/DRAM_ADDR_net_0[15] , 
        \SF2Project_MSS_0/DRAM_ADDR_net_0[14] , 
        \SF2Project_MSS_0/DRAM_ADDR_net_0[13] , 
        \SF2Project_MSS_0/DRAM_ADDR_net_0[12] , 
        \SF2Project_MSS_0/DRAM_ADDR_net_0[11] , 
        \SF2Project_MSS_0/DRAM_ADDR_net_0[10] , 
        \SF2Project_MSS_0/DRAM_ADDR_net_0[9] , 
        \SF2Project_MSS_0/DRAM_ADDR_net_0[8] , 
        \SF2Project_MSS_0/DRAM_ADDR_net_0[7] , 
        \SF2Project_MSS_0/DRAM_ADDR_net_0[6] , 
        \SF2Project_MSS_0/DRAM_ADDR_net_0[5] , 
        \SF2Project_MSS_0/DRAM_ADDR_net_0[4] , 
        \SF2Project_MSS_0/DRAM_ADDR_net_0[3] , 
        \SF2Project_MSS_0/DRAM_ADDR_net_0[2] , 
        \SF2Project_MSS_0/DRAM_ADDR_net_0[1] , 
        \SF2Project_MSS_0/DRAM_ADDR_net_0[0] , 
        \SF2Project_MSS_0/DRAM_DQS_OUT_net_0[1] , 
        \SF2Project_MSS_0/DRAM_DQS_OUT_net_0[0] , 
        \SF2Project_MSS_0/DRAM_DQS_OE_net_0[1] , 
        \SF2Project_MSS_0/DRAM_DQS_OE_net_0[0] , 
        \SF2Project_MSS_0/USB_ULPI_XCLK_PAD_Y , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_TXD1_RMII_TXD1_USBB_STP_OUT , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_TXD1_RMII_TXD1_USBB_STP_OE , 
        \SF2Project_MSS_0/USB_ULPI_NXT_PAD_Y , 
        \SF2Project_MSS_0/USB_ULPI_DIR_PAD_Y , 
        \SF2Project_MSS_0/USB_ULPI_DATA_7_PAD_Y , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE , 
        \SF2Project_MSS_0/USB_ULPI_DATA_6_PAD_Y , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_TXD3_USBB_DATA6_OUT , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_TXD3_USBB_DATA6_OE , 
        \SF2Project_MSS_0/USB_ULPI_DATA_5_PAD_Y , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_TXD2_USBB_DATA5_OUT , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_TXD2_USBB_DATA5_OE , 
        \SF2Project_MSS_0/USB_ULPI_DATA_4_PAD_Y , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_RXD3_USBB_DATA4_OUT , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_RXD3_USBB_DATA4_OE , 
        \SF2Project_MSS_0/USB_ULPI_DATA_3_PAD_Y , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE , 
        \SF2Project_MSS_0/USB_ULPI_DATA_2_PAD_Y , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE , 
        \SF2Project_MSS_0/USB_ULPI_DATA_1_PAD_Y , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE , 
        \SF2Project_MSS_0/USB_ULPI_DATA_0_PAD_Y , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE , 
        \SF2Project_MSS_0/SPI_1_SS0_PAD_Y , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_SPI1_SS0_MGPIO13A_OUT , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_SPI1_SS0_MGPIO13A_OE , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_SPI1_SDO_MGPIO12A_OUT , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_SPI1_SDO_MGPIO12A_OE , 
        \SF2Project_MSS_0/SPI_1_DI_PAD_Y , 
        \SF2Project_MSS_0/SPI_1_CLK_PAD_Y , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_SPI1_SCK_OUT , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_SPI1_SCK_OE , 
        \SF2Project_MSS_0/SPI_0_SS0_PAD_Y , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OUT , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OE , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OUT , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OE , 
        \SF2Project_MSS_0/SPI_0_DI_PAD_Y , 
        \SF2Project_MSS_0/SPI_0_CLK_PAD_Y , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OUT , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OE , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OE , 
        \SF2Project_MSS_0/MMUART_1_RXD_PAD_Y , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OUT , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OE , 
        \SF2Project_MSS_0/MMUART_0_RXD_PAD_Y , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_DRAM_WEN , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_DRAM_RSTN , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_DRAM_RASN , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_DRAM_ODT , 
        \SF2Project_MSS_0/MDDR_DQS_TMATCH_0_IN_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DQ_15_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DQ_14_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DQ_13_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DQ_12_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DQ_11_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DQ_10_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DQ_9_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DQ_8_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DQ_7_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DQ_6_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DQ_5_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DQ_4_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DQ_3_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DQ_2_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DQ_1_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DQ_0_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DM_RDQS_1_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DM_RDQS_0_PAD_Y , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_DRAM_CSN , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_DRAM_CKE , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_DRAM_CASN , 
        \SF2Project_MSS_0/I2C_1_SDA_PAD_Y , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OUT , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OE , 
        \SF2Project_MSS_0/I2C_1_SCL_PAD_Y , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OUT , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OE , 
        \SF2Project_MSS_0/I2C_0_SDA_PAD_Y , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_I2C0_SDA_USBC_DATA0_MGPIO30B_OUT , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_I2C0_SDA_USBC_DATA0_MGPIO30B_OE , 
        \SF2Project_MSS_0/I2C_0_SCL_PAD_Y , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_I2C0_SCL_USBC_DATA1_MGPIO31B_OUT , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_I2C0_SCL_USBC_DATA1_MGPIO31B_OE , 
        VCC, GND, \SF2Project_MSS_0/MDDR_DQS_0_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DQS_1_PAD_Y , 
        \SF2Project_MSS_0/MSS_ADLIB_INST_DRAM_CLK , 
        \SF2Project_MSS_0/MDDR_ODT_PAD/EOUT , 
        \SF2Project_MSS_0/MDDR_BA_0_PAD/EOUT , 
        \SF2Project_MSS_0/MDDR_WE_N_PAD/EOUT , 
        \SF2Project_MSS_0/USB_ULPI_DATA_7_PAD/YIN , 
        \SF2Project_MSS_0/USB_ULPI_DATA_0_PAD/YIN , 
        \SF2Project_MSS_0/MDDR_RESET_N_PAD/EOUT , 
        \SF2Project_MSS_0/SPI_0_SS0_PAD/YIN , 
        \SF2Project_MSS_0/MDDR_DM_RDQS_1_PAD/YIN , 
        \SF2Project_MSS_0/MDDR_ADDR_9_PAD/EOUT , 
        \SF2Project_MSS_0/MDDR_DQ_4_PAD/YIN , 
        \SF2Project_MSS_0/SPI_1_DI_PAD/YIN , 
        \SF2Project_MSS_0/MMUART_0_RXD_PAD/YIN , 
        \SF2Project_MSS_0/MMUART_1_RXD_PAD/YIN , 
        \SF2Project_MSS_0/MDDR_DQ_5_PAD/YIN , 
        \SF2Project_MSS_0/USB_ULPI_DIR_PAD/YIN , 
        \SF2Project_MSS_0/MDDR_ADDR_0_PAD/EOUT , 
        \SF2Project_MSS_0/USB_ULPI_NXT_PAD/YIN , 
        \SF2Project_MSS_0/MDDR_DQ_9_PAD/YIN , 
        \SF2Project_MSS_0/SPI_1_SS0_PAD/YIN , 
        \SF2Project_MSS_0/SPI_0_CLK_PAD/YIN , 
        \SF2Project_MSS_0/MDDR_DQ_1_PAD/YIN , 
        \SF2Project_MSS_0/MDDR_ADDR_2_PAD/EOUT , 
        \SF2Project_MSS_0/MDDR_BA_1_PAD/EOUT , 
        \SF2Project_MSS_0/MDDR_ADDR_6_PAD/EOUT , 
        \SF2Project_MSS_0/MDDR_DQ_7_PAD/YIN , 
        \SF2Project_MSS_0/MDDR_ADDR_4_PAD/EOUT , 
        \SF2Project_MSS_0/MDDR_DQ_2_PAD/YIN , 
        \SF2Project_MSS_0/MDDR_ADDR_1_PAD/EOUT , 
        \SF2Project_MSS_0/MDDR_DQS_1_PAD/U2_N2P , 
        \SF2Project_MSS_0/MDDR_DQS_1_PAD/YIN , 
        \SF2Project_MSS_0/MDDR_ADDR_15_PAD/EOUT , 
        \SF2Project_MSS_0/MDDR_CS_N_PAD/EOUT , 
        \SF2Project_MSS_0/MDDR_ADDR_8_PAD/EOUT , 
        \SF2Project_MSS_0/USB_ULPI_XCLK_PAD/YIN , 
        \SF2Project_MSS_0/MDDR_DQ_11_PAD/YIN , 
        \SF2Project_MSS_0/MDDR_ADDR_10_PAD/EOUT , 
        \SF2Project_MSS_0/MDDR_DQS_0_PAD/U2_N2P , 
        \SF2Project_MSS_0/MDDR_DQS_0_PAD/YIN , 
        \SF2Project_MSS_0/MDDR_CAS_N_PAD/EOUT , 
        \SF2Project_MSS_0/MDDR_BA_2_PAD/EOUT , 
        \SF2Project_MSS_0/USB_ULPI_DATA_4_PAD/YIN , 
        \SF2Project_MSS_0/I2C_1_SCL_PAD/YIN , 
        \SF2Project_MSS_0/USB_ULPI_DATA_2_PAD/YIN , 
        \SF2Project_MSS_0/USB_ULPI_DATA_3_PAD/YIN , 
        \SF2Project_MSS_0/MDDR_RAS_N_PAD/EOUT , 
        \SF2Project_MSS_0/MDDR_DQS_TMATCH_0_IN_PAD/YIN , 
        \SF2Project_MSS_0/MDDR_DQ_8_PAD/YIN , 
        \SF2Project_MSS_0/MDDR_ADDR_5_PAD/EOUT , 
        \SF2Project_MSS_0/MDDR_DQ_15_PAD/YIN , 
        \SF2Project_MSS_0/I2C_1_SDA_PAD/YIN , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/CAN_RXBUS_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/CAN_TX_EBL_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/CAN_TXBUS_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/COLF_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/CRSF_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2_DMAREADY_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2_DMAREADY_net[0] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[15] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[14] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[13] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[12] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[11] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[10] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[9] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[8] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[7] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[6] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[5] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[4] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[0] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2HCALIB_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_DMAREADY_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_DMAREADY_net[0] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[31] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[30] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[29] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[28] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[27] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[26] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[25] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[24] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[23] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[22] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[21] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[20] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[19] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[18] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[17] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[16] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[15] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[14] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[13] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[12] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[11] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[10] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[9] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[8] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[7] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[6] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[5] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[4] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[0] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ENABLE_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_MASTLOCK_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_READY_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_SEL_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_SIZE_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_SIZE_net[0] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_TRANS1_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[31] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[30] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[29] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[28] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[27] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[26] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[25] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[24] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[23] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[22] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[21] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[20] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[19] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[18] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[17] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[16] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[15] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[14] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[13] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[12] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[11] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[10] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[9] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[8] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[7] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[6] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[5] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[4] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[0] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WRITE_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[31] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[30] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[29] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[28] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[27] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[26] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[25] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[24] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[23] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[22] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[21] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[20] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[19] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[18] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[17] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[16] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[15] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[14] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[13] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[12] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[11] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[10] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[9] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[8] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[7] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[6] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[5] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[4] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[0] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_READY_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RESP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_AVALID_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_HOSTDISCON_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_IDDIG_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_LINESTATE_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_LINESTATE_net[0] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_M3_RESET_N_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_PLL_LOCK_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_RXACTIVE_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_RXERROR_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_RXVALID_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_RXVALIDH_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_SESSEND_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_TXREADY_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_VBUSVALID_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[7] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[6] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[5] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[4] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[0] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[7] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[6] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[5] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[4] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[0] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/GTX_CLKPF_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/I2C0_BCLK_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/I2C0_SCL_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/I2C0_SDA_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/I2C1_BCLK_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/I2C1_SCL_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/I2C1_SDA_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDIF_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO0A_F2H_GPIN_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO10A_F2H_GPIN_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO11A_F2H_GPIN_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO11B_F2H_GPIN_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO12A_F2H_GPIN_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO13A_F2H_GPIN_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO14A_F2H_GPIN_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO15A_F2H_GPIN_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO16A_F2H_GPIN_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO17B_F2H_GPIN_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO18B_F2H_GPIN_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO19B_F2H_GPIN_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO1A_F2H_GPIN_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO20B_F2H_GPIN_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO21B_F2H_GPIN_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO22B_F2H_GPIN_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO24B_F2H_GPIN_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO25B_F2H_GPIN_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO26B_F2H_GPIN_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO27B_F2H_GPIN_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO28B_F2H_GPIN_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO29B_F2H_GPIN_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO2A_F2H_GPIN_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO30B_F2H_GPIN_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO31B_F2H_GPIN_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO3A_F2H_GPIN_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO4A_F2H_GPIN_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO5A_F2H_GPIN_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO6A_F2H_GPIN_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO7A_F2H_GPIN_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO8A_F2H_GPIN_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO9A_F2H_GPIN_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART0_CTS_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART0_DCD_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART0_DSR_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART0_DTR_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART0_RI_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART0_RTS_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART0_RXD_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART0_SCK_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART0_TXD_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART1_CTS_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART1_DCD_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART1_DSR_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART1_RI_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART1_RTS_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART1_RXD_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART1_SCK_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART1_TXD_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[31] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[30] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[29] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[28] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[27] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[26] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[25] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[24] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[23] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[22] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[21] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[20] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[19] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[18] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[17] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[16] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[15] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[14] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[13] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[12] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[11] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[10] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[9] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[8] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[7] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[6] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[5] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[4] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[0] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PREADY_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PSLVERR_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RCGF_net[9] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RCGF_net[8] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RCGF_net[7] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RCGF_net[6] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RCGF_net[5] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RCGF_net[4] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RCGF_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RCGF_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RCGF_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RCGF_net[0] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RX_CLKPF_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RX_DVF_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RX_ERRF_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RX_EV_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RXDF_net[7] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RXDF_net[6] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RXDF_net[5] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RXDF_net[4] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RXDF_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RXDF_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RXDF_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RXDF_net[0] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/SLEEPHOLDREQ_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/SMBALERT_NI0_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/SMBALERT_NI1_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/SMBSUS_NI0_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/SMBSUS_NI1_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI0_CLK_IN_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI0_SDI_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI0_SDO_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI0_SS0_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI0_SS1_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI0_SS2_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI0_SS3_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI1_CLK_IN_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI1_SDI_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI1_SDO_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI1_SS0_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI1_SS1_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI1_SS2_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI1_SS3_F2H_SCP_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/TX_CLKPF_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/USER_MSS_GPIO_RESET_N_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/USER_MSS_RESET_N_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/XCLK_FAB_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/CLK_BASE_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/CLK_MDDR_APB_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[31] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[30] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[29] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[28] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[27] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[26] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[25] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[24] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[23] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[22] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[21] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[20] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[19] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[18] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[17] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[16] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[15] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[14] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[13] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[12] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[11] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[10] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[9] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[8] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[7] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[6] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[5] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[4] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[0] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARBURST_HTRANS1_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARBURST_HTRANS1_net[0] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[0] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[0] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARLOCK_HMASTLOCK1_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARLOCK_HMASTLOCK1_net[0] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARSIZE_HSIZE1_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARSIZE_HSIZE1_net[0] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARVALID_HWRITE1_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[31] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[30] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[29] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[28] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[27] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[26] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[25] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[24] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[23] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[22] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[21] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[20] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[19] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[18] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[17] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[16] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[15] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[14] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[13] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[12] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[11] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[10] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[9] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[8] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[7] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[6] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[5] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[4] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[0] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWBURST_HTRANS0_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWBURST_HTRANS0_net[0] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[0] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[0] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWLOCK_HMASTLOCK0_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWLOCK_HMASTLOCK0_net[0] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWSIZE_HSIZE0_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWSIZE_HSIZE0_net[0] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWVALID_HWRITE0_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_BREADY_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_RMW_AXI_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_RREADY_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[63] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[62] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[61] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[60] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[59] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[58] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[57] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[56] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[55] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[54] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[53] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[52] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[51] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[50] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[49] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[48] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[47] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[46] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[45] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[44] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[43] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[42] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[41] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[40] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[39] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[38] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[37] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[36] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[35] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[34] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[33] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[32] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[31] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[30] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[29] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[28] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[27] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[26] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[25] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[24] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[23] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[22] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[21] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[20] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[19] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[18] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[17] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[16] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[15] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[14] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[13] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[12] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[11] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[10] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[9] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[8] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[7] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[6] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[5] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[4] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[0] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[0] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WLAST_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[7] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[6] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[5] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[4] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[0] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WVALID_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FPGA_MDDR_ARESET_N_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[10] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[9] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[8] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[7] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[6] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[5] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[4] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PENABLE_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PSEL_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[15] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[14] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[13] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[12] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[11] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[10] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[9] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[8] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[7] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[6] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[5] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[4] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[0] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWRITE_net , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PRESET_N_net , 
        \SF2Project_MSS_0/MDDR_DQ_0_PAD/YIN , 
        \SF2Project_MSS_0/MDDR_ADDR_13_PAD/EOUT , 
        \SF2Project_MSS_0/MDDR_DM_RDQS_0_PAD/YIN , 
        \SF2Project_MSS_0/MDDR_ADDR_14_PAD/EOUT , 
        \SF2Project_MSS_0/MDDR_DQ_13_PAD/YIN , 
        \SF2Project_MSS_0/MDDR_ADDR_12_PAD/EOUT , 
        \SF2Project_MSS_0/MDDR_DQ_14_PAD/YIN , 
        \SF2Project_MSS_0/MDDR_DQ_6_PAD/YIN , 
        \SF2Project_MSS_0/USB_ULPI_DATA_5_PAD/YIN , 
        \SF2Project_MSS_0/MDDR_ADDR_7_PAD/EOUT , 
        \SF2Project_MSS_0/MDDR_ADDR_11_PAD/EOUT , 
        \SF2Project_MSS_0/USB_ULPI_DATA_1_PAD/YIN , 
        \SF2Project_MSS_0/MDDR_CKE_PAD/EOUT , 
        \SF2Project_MSS_0/I2C_0_SDA_PAD/YIN , 
        \SF2Project_MSS_0/USB_ULPI_DATA_6_PAD/YIN , 
        \SF2Project_MSS_0/SPI_0_DI_PAD/YIN , 
        \SF2Project_MSS_0/MDDR_DQ_12_PAD/YIN , 
        \SF2Project_MSS_0/SPI_1_CLK_PAD/YIN , 
        \SF2Project_MSS_0/MDDR_DQ_3_PAD/YIN , 
        \SF2Project_MSS_0/I2C_0_SCL_PAD/YIN , 
        \SF2Project_MSS_0/MDDR_DQS_TMATCH_0_OUT_PAD/EOUT , 
        \SF2Project_MSS_0/MDDR_ADDR_3_PAD/EOUT , 
        \SF2Project_MSS_0/MDDR_DQ_10_PAD/YIN , AFLSDF_VCC, AFLSDF_GND;
    wire GND_power_net1;
    wire VCC_power_net1;
    assign GND = GND_power_net1;
    assign AFLSDF_GND = GND_power_net1;
    assign VCC = VCC_power_net1;
    assign AFLSDF_VCC = VCC_power_net1;
    
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_17  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[22] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[29] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_110  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[2] ), .IPB(), 
        .IPC());
    IOIN_IB \SF2Project_MSS_0/USB_ULPI_DIR_PAD/U_IOIN  (.YIN(
        \SF2Project_MSS_0/USB_ULPI_DIR_PAD/YIN ), .E(GND), .Y());
    sdf_IOPAD_TRI \SF2Project_MSS_0/MDDR_ADDR_1_PAD/U_IOPAD  (.PAD(
        MDDR_ADDR[1]), .D(\SF2Project_MSS_0/DRAM_ADDR_net_0[1] ), .E(
        \SF2Project_MSS_0/MDDR_ADDR_1_PAD/EOUT ));
    IOBI_IB_OB_EB \SF2Project_MSS_0/MDDR_DQ_5_PAD/U_IOBI  (.D(VCC), .E(
        VCC), .YIN(\SF2Project_MSS_0/MDDR_DQ_5_PAD/YIN ), .DOUT(), 
        .EOUT(), .Y());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_85  (.A(
        VCC), .B(\MAC_MII_RXD[1] ), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[26] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/RXDF_net[1] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_64  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[25] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PREADY_net ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_81  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[15] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[22] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_40  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[23] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[30] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_182  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO27B_F2H_GPIN_net ), .IPB(
        ), .IPC());
    IOBI_IB_OB_EB \SF2Project_MSS_0/MDDR_DQ_6_PAD/U_IOBI  (.D(VCC), .E(
        VCC), .YIN(\SF2Project_MSS_0/MDDR_DQ_6_PAD/YIN ), .DOUT(), 
        .EOUT(), .Y());
    IOTRI_OB_EB \SF2Project_MSS_0/MDDR_ADDR_13_PAD/U_IOOUT  (.D(VCC), 
        .E(VCC), .DOUT(), .EOUT(
        \SF2Project_MSS_0/MDDR_ADDR_13_PAD/EOUT ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_269  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[29] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_ARVALID_HWRITE1_net ), 
        .IPC());
    IOINFF_BYPASS \SF2Project_MSS_0/USB_ULPI_DATA_7_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/USB_ULPI_DATA_7_PAD_Y ), .Y(
        \SF2Project_MSS_0/USB_ULPI_DATA_7_PAD/YIN ));
    sdf_IOPAD_TRI \SF2Project_MSS_0/SPI_1_DO_PAD/U_IOPAD  (.PAD(
        SPI_1_DO), .D(
        \SF2Project_MSS_0/MSS_ADLIB_INST_SPI1_SDO_MGPIO12A_OUT ), .E(
        \SF2Project_MSS_0/MSS_ADLIB_INST_SPI1_SDO_MGPIO12A_OE ));
    sdf_IOPAD_TRI \SF2Project_MSS_0/MDDR_CAS_N_PAD/U_IOPAD  (.PAD(
        MDDR_CAS_N), .D(\SF2Project_MSS_0/MSS_ADLIB_INST_DRAM_CASN ), 
        .E(\SF2Project_MSS_0/MDDR_CAS_N_PAD/EOUT ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_98  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDIF_net ), .IPB(), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_274  (
        .A(GND), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[2] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/CLK_MDDR_APB_net ), .IPC(
        ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_174  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO25B_F2H_GPIN_net ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART0_DTR_F2H_SCP_net ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_16  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[21] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[28] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_57  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[11] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[18] ), .IPC());
    sdf_IOPAD_TRI \SF2Project_MSS_0/MDDR_ADDR_9_PAD/U_IOPAD  (.PAD(
        MDDR_ADDR[9]), .D(\SF2Project_MSS_0/DRAM_ADDR_net_0[9] ), .E(
        \SF2Project_MSS_0/MDDR_ADDR_9_PAD/EOUT ));
    IOTRI_OB_EB \SF2Project_MSS_0/MDDR_ADDR_9_PAD/U_IOOUT  (.D(VCC), 
        .E(VCC), .DOUT(), .EOUT(
        \SF2Project_MSS_0/MDDR_ADDR_9_PAD/EOUT ));
    sdf_IOPADN_BI \SF2Project_MSS_0/MDDR_DQS_0_PAD/U_IOPADN  (.PAD_P(
        MDDR_DQS_N[0]), .OIN_P(
        \SF2Project_MSS_0/DRAM_DQS_OUT_net_0[0] ), .EIN_P(
        \SF2Project_MSS_0/DRAM_DQS_OE_net_0[0] ), .N2POUT_P(
        \SF2Project_MSS_0/MDDR_DQS_0_PAD/U2_N2P ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_179  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO21B_F2H_GPIN_net ), .IPC(
        ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_68  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[29] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[2] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_37  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[20] ), .IPB(), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_105  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/RCGF_net[5] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_LINESTATE_net[1] ), .IPC()
        );
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_170  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART1_RI_F2H_SCP_net ), 
        .IPB(), .IPC());
    IOTRI_OB_EB \SF2Project_MSS_0/MDDR_BA_1_PAD/U_IOOUT  (.D(VCC), .E(
        VCC), .DOUT(), .EOUT(\SF2Project_MSS_0/MDDR_BA_1_PAD/EOUT ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_264  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[24] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARBURST_HTRANS1_net[0] ), 
        .IPC(\SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PENABLE_net )
        );
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_164  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO13A_F2H_GPIN_net ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO16A_F2H_GPIN_net ), .IPC(
        ));
    IOBI_IB_OB_EB \SF2Project_MSS_0/SPI_1_SS0_PAD/U_IOBI  (.D(VCC), .E(
        VCC), .YIN(\SF2Project_MSS_0/SPI_1_SS0_PAD/YIN ), .DOUT(), 
        .EOUT(), .Y());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_56  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[10] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[17] ), .IPC());
    MSS_010_IP #( .INIT(1438'h0000040100361200000000000000003610008000000000000000000000000000000000001203610000000000000000000120361000000000100520481204812048120D8120D8120F00000000F000000000000000000000000000000007FFFFFFFB000001007C37F00020200E09280F00183FFFFE400000000002150000000000E11C0000007E4800010842108421000001FE34001FF8000000400000000020091007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
        , .ACT_UBITS(56'hFFFFFFFFFFFFFF), .MEMORYFILE("ENVM_init.mem")
        , .RTC_MAIN_XTL_FREQ(0.000000), .RTC_MAIN_XTL_MODE(""), .DDR_CLK_FREQ(200.000000)
         )  \SF2Project_MSS_0/MSS_ADLIB_INST/INST_MSS_010_IP  (
        .CAN_RXBUS_MGPIO3A_H2F_A(), .CAN_RXBUS_MGPIO3A_H2F_B(), 
        .CAN_TX_EBL_MGPIO4A_H2F_A(), .CAN_TX_EBL_MGPIO4A_H2F_B(), 
        .CAN_TXBUS_MGPIO2A_H2F_A(), .CAN_TXBUS_MGPIO2A_H2F_B(), 
        .CLK_CONFIG_APB(), .COMMS_INT(), .CONFIG_PRESET_N(), 
        .EDAC_ERROR({nc0, nc1, nc2, nc3, nc4, nc5, nc6, nc7}), 
        .F_FM0_RDATA({nc8, nc9, nc10, nc11, nc12, nc13, nc14, nc15, 
        nc16, nc17, nc18, nc19, nc20, nc21, nc22, nc23, nc24, nc25, 
        nc26, nc27, nc28, nc29, nc30, nc31, nc32, nc33, nc34, nc35, 
        nc36, nc37, nc38, nc39}), .F_FM0_READYOUT(), .F_FM0_RESP(), 
        .F_HM0_ADDR({nc40, nc41, nc42, nc43, nc44, nc45, nc46, nc47, 
        nc48, nc49, nc50, nc51, nc52, nc53, nc54, nc55, nc56, nc57, 
        nc58, nc59, nc60, nc61, nc62, nc63, nc64, nc65, nc66, nc67, 
        nc68, nc69, nc70, nc71}), .F_HM0_ENABLE(), .F_HM0_SEL(), 
        .F_HM0_SIZE({nc72, nc73}), .F_HM0_TRANS1(), .F_HM0_WDATA({nc74, 
        nc75, nc76, nc77, nc78, nc79, nc80, nc81, nc82, nc83, nc84, 
        nc85, nc86, nc87, nc88, nc89, nc90, nc91, nc92, nc93, nc94, 
        nc95, nc96, nc97, nc98, nc99, nc100, nc101, nc102, nc103, 
        nc104, nc105}), .F_HM0_WRITE(), .FAB_CHRGVBUS(), 
        .FAB_DISCHRGVBUS(), .FAB_DMPULLDOWN(), .FAB_DPPULLDOWN(), 
        .FAB_DRVVBUS(), .FAB_IDPULLUP(), .FAB_OPMODE({nc106, nc107}), 
        .FAB_SUSPENDM(), .FAB_TERMSEL(), .FAB_TXVALID(), .FAB_VCONTROL({
        nc108, nc109, nc110, nc111}), .FAB_VCONTROLLOADM(), 
        .FAB_XCVRSEL({nc112, nc113}), .FAB_XDATAOUT({nc114, nc115, 
        nc116, nc117, nc118, nc119, nc120, nc121}), .FACC_GLMUX_SEL(), 
        .FIC32_0_MASTER({nc122, nc123}), .FIC32_1_MASTER({nc124, nc125})
        , .FPGA_RESET_N(), .GTX_CLK(), .H2F_INTERRUPT({nc126, nc127, 
        nc128, nc129, nc130, nc131, nc132, nc133, nc134, nc135, nc136, 
        nc137, nc138, nc139, nc140, nc141}), .H2F_NMI(), .H2FCALIB(), 
        .I2C0_SCL_MGPIO31B_H2F_A(), .I2C0_SCL_MGPIO31B_H2F_B(), 
        .I2C0_SDA_MGPIO30B_H2F_A(), .I2C0_SDA_MGPIO30B_H2F_B(), 
        .I2C1_SCL_MGPIO1A_H2F_A(), .I2C1_SCL_MGPIO1A_H2F_B(), 
        .I2C1_SDA_MGPIO0A_H2F_A(), .I2C1_SDA_MGPIO0A_H2F_B(), .MDCF(), 
        .MDOENF(), .MDOF(), .MMUART0_CTS_MGPIO19B_H2F_A(), 
        .MMUART0_CTS_MGPIO19B_H2F_B(), .MMUART0_DCD_MGPIO22B_H2F_A(), 
        .MMUART0_DCD_MGPIO22B_H2F_B(), .MMUART0_DSR_MGPIO20B_H2F_A(), 
        .MMUART0_DSR_MGPIO20B_H2F_B(), .MMUART0_DTR_MGPIO18B_H2F_A(), 
        .MMUART0_DTR_MGPIO18B_H2F_B(), .MMUART0_RI_MGPIO21B_H2F_A(), 
        .MMUART0_RI_MGPIO21B_H2F_B(), .MMUART0_RTS_MGPIO17B_H2F_A(), 
        .MMUART0_RTS_MGPIO17B_H2F_B(), .MMUART0_RXD_MGPIO28B_H2F_A(), 
        .MMUART0_RXD_MGPIO28B_H2F_B(), .MMUART0_SCK_MGPIO29B_H2F_A(), 
        .MMUART0_SCK_MGPIO29B_H2F_B(), .MMUART0_TXD_MGPIO27B_H2F_A(), 
        .MMUART0_TXD_MGPIO27B_H2F_B(), .MMUART1_DTR_MGPIO12B_H2F_A(), 
        .MMUART1_RTS_MGPIO11B_H2F_A(), .MMUART1_RTS_MGPIO11B_H2F_B(), 
        .MMUART1_RXD_MGPIO26B_H2F_A(), .MMUART1_RXD_MGPIO26B_H2F_B(), 
        .MMUART1_SCK_MGPIO25B_H2F_A(), .MMUART1_SCK_MGPIO25B_H2F_B(), 
        .MMUART1_TXD_MGPIO24B_H2F_A(), .MMUART1_TXD_MGPIO24B_H2F_B(), 
        .MPLL_LOCK(), .PER2_FABRIC_PADDR({nc142, nc143, nc144, nc145, 
        nc146, nc147, nc148, nc149, nc150, nc151, nc152, nc153, nc154, 
        nc155}), .PER2_FABRIC_PENABLE(), .PER2_FABRIC_PSEL(), 
        .PER2_FABRIC_PWDATA({nc156, nc157, nc158, nc159, nc160, nc161, 
        nc162, nc163, nc164, nc165, nc166, nc167, nc168, nc169, nc170, 
        nc171, nc172, nc173, nc174, nc175, nc176, nc177, nc178, nc179, 
        nc180, nc181, nc182, nc183, nc184, nc185, nc186, nc187}), 
        .PER2_FABRIC_PWRITE(), .RTC_MATCH(), .SLEEPDEEP(), 
        .SLEEPHOLDACK(), .SLEEPING(), .SMBALERT_NO0(), .SMBALERT_NO1(), 
        .SMBSUS_NO0(), .SMBSUS_NO1(), .SPI0_CLK_OUT(), 
        .SPI0_SDI_MGPIO5A_H2F_A(), .SPI0_SDI_MGPIO5A_H2F_B(), 
        .SPI0_SDO_MGPIO6A_H2F_A(), .SPI0_SDO_MGPIO6A_H2F_B(), 
        .SPI0_SS0_MGPIO7A_H2F_A(), .SPI0_SS0_MGPIO7A_H2F_B(), 
        .SPI0_SS1_MGPIO8A_H2F_A(), .SPI0_SS1_MGPIO8A_H2F_B(), 
        .SPI0_SS2_MGPIO9A_H2F_A(), .SPI0_SS2_MGPIO9A_H2F_B(), 
        .SPI0_SS3_MGPIO10A_H2F_A(), .SPI0_SS3_MGPIO10A_H2F_B(), 
        .SPI0_SS4_MGPIO19A_H2F_A(), .SPI0_SS5_MGPIO20A_H2F_A(), 
        .SPI0_SS6_MGPIO21A_H2F_A(), .SPI0_SS7_MGPIO22A_H2F_A(), 
        .SPI1_CLK_OUT(), .SPI1_SDI_MGPIO11A_H2F_A(), 
        .SPI1_SDI_MGPIO11A_H2F_B(), .SPI1_SDO_MGPIO12A_H2F_A(), 
        .SPI1_SDO_MGPIO12A_H2F_B(), .SPI1_SS0_MGPIO13A_H2F_A(), 
        .SPI1_SS0_MGPIO13A_H2F_B(), .SPI1_SS1_MGPIO14A_H2F_A(), 
        .SPI1_SS1_MGPIO14A_H2F_B(), .SPI1_SS2_MGPIO15A_H2F_A(), 
        .SPI1_SS2_MGPIO15A_H2F_B(), .SPI1_SS3_MGPIO16A_H2F_A(), 
        .SPI1_SS3_MGPIO16A_H2F_B(), .SPI1_SS4_MGPIO17A_H2F_A(), 
        .SPI1_SS5_MGPIO18A_H2F_A(), .SPI1_SS6_MGPIO23A_H2F_A(), 
        .SPI1_SS7_MGPIO24A_H2F_A(), .TCGF({nc188, nc189, nc190, nc191, 
        nc192, nc193, nc194, nc195, nc196, nc197}), .TRACECLK(), 
        .TRACEDATA({nc198, nc199, nc200, nc201}), .TX_CLK(), .TX_ENF(
        MAC_MII_TX_EN_net_1), .TX_ERRF(MAC_MII_TX_ER_net_1), 
        .TXCTL_EN_RIF(), .TXD_RIF({nc202, nc203, nc204, nc205}), .TXDF({
        nc206, nc207, nc208, nc209, \MAC_MII_TXD[3] , \MAC_MII_TXD[2] , 
        \MAC_MII_TXD[1] , \MAC_MII_TXD[0] }), .TXEV(), .WDOGTIMEOUT(), 
        .F_ARREADY_HREADYOUT1(), .F_AWREADY_HREADYOUT0(), .F_BID({
        nc210, nc211, nc212, nc213}), .F_BRESP_HRESP0({nc214, nc215}), 
        .F_BVALID(), .F_RDATA_HRDATA01({nc216, nc217, nc218, nc219, 
        nc220, nc221, nc222, nc223, nc224, nc225, nc226, nc227, nc228, 
        nc229, nc230, nc231, nc232, nc233, nc234, nc235, nc236, nc237, 
        nc238, nc239, nc240, nc241, nc242, nc243, nc244, nc245, nc246, 
        nc247, nc248, nc249, nc250, nc251, nc252, nc253, nc254, nc255, 
        nc256, nc257, nc258, nc259, nc260, nc261, nc262, nc263, nc264, 
        nc265, nc266, nc267, nc268, nc269, nc270, nc271, nc272, nc273, 
        nc274, nc275, nc276, nc277, nc278, nc279}), .F_RID({nc280, 
        nc281, nc282, nc283}), .F_RLAST(), .F_RRESP_HRESP1({nc284, 
        nc285}), .F_RVALID(), .F_WREADY(), .MDDR_FABRIC_PRDATA({nc286, 
        nc287, nc288, nc289, nc290, nc291, nc292, nc293, nc294, nc295, 
        nc296, nc297, nc298, nc299, nc300, nc301}), 
        .MDDR_FABRIC_PREADY(), .MDDR_FABRIC_PSLVERR(), 
        .CAN_RXBUS_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/CAN_RXBUS_F2H_SCP_net ), 
        .CAN_TX_EBL_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/CAN_TX_EBL_F2H_SCP_net ), 
        .CAN_TXBUS_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/CAN_TXBUS_F2H_SCP_net ), 
        .COLF(\SF2Project_MSS_0/MSS_ADLIB_INST/COLF_net ), .CRSF(
        \SF2Project_MSS_0/MSS_ADLIB_INST/CRSF_net ), .F2_DMAREADY({
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2_DMAREADY_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2_DMAREADY_net[0] }), 
        .F2H_INTERRUPT({
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[15] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[14] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[13] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[12] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[11] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[10] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[9] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[8] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[7] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[6] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[5] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[4] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[0] }), 
        .F2HCALIB(\SF2Project_MSS_0/MSS_ADLIB_INST/F2HCALIB_net ), 
        .F_DMAREADY({
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_DMAREADY_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_DMAREADY_net[0] }), 
        .F_FM0_ADDR({
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[31] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[30] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[29] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[28] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[27] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[26] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[25] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[24] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[23] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[22] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[21] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[20] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[19] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[18] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[17] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[16] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[15] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[14] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[13] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[12] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[11] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[10] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[9] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[8] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[7] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[6] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[5] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[4] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[0] }), 
        .F_FM0_ENABLE(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ENABLE_net ), 
        .F_FM0_MASTLOCK(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_MASTLOCK_net ), 
        .F_FM0_READY(\SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_READY_net )
        , .F_FM0_SEL(\SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_SEL_net ), 
        .F_FM0_SIZE({
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_SIZE_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_SIZE_net[0] }), 
        .F_FM0_TRANS1(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_TRANS1_net ), 
        .F_FM0_WDATA({
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[31] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[30] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[29] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[28] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[27] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[26] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[25] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[24] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[23] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[22] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[21] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[20] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[19] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[18] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[17] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[16] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[15] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[14] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[13] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[12] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[11] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[10] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[9] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[8] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[7] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[6] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[5] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[4] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[0] }), 
        .F_FM0_WRITE(\SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WRITE_net )
        , .F_HM0_RDATA({
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[31] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[30] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[29] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[28] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[27] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[26] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[25] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[24] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[23] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[22] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[21] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[20] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[19] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[18] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[17] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[16] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[15] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[14] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[13] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[12] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[11] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[10] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[9] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[8] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[7] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[6] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[5] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[4] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[0] }), 
        .F_HM0_READY(\SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_READY_net )
        , .F_HM0_RESP(\SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RESP_net )
        , .FAB_AVALID(\SF2Project_MSS_0/MSS_ADLIB_INST/FAB_AVALID_net )
        , .FAB_HOSTDISCON(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_HOSTDISCON_net ), 
        .FAB_IDDIG(\SF2Project_MSS_0/MSS_ADLIB_INST/FAB_IDDIG_net ), 
        .FAB_LINESTATE({
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_LINESTATE_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_LINESTATE_net[0] }), 
        .FAB_M3_RESET_N(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_M3_RESET_N_net ), 
        .FAB_PLL_LOCK(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_PLL_LOCK_net ), 
        .FAB_RXACTIVE(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_RXACTIVE_net ), 
        .FAB_RXERROR(\SF2Project_MSS_0/MSS_ADLIB_INST/FAB_RXERROR_net )
        , .FAB_RXVALID(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_RXVALID_net ), 
        .FAB_RXVALIDH(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_RXVALIDH_net ), 
        .FAB_SESSEND(\SF2Project_MSS_0/MSS_ADLIB_INST/FAB_SESSEND_net )
        , .FAB_TXREADY(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_TXREADY_net ), 
        .FAB_VBUSVALID(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_VBUSVALID_net ), 
        .FAB_VSTATUS({
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[7] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[6] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[5] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[4] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[0] }), 
        .FAB_XDATAIN({
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[7] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[6] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[5] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[4] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[0] }), 
        .GTX_CLKPF(\SF2Project_MSS_0/MSS_ADLIB_INST/GTX_CLKPF_net ), 
        .I2C0_BCLK(\SF2Project_MSS_0/MSS_ADLIB_INST/I2C0_BCLK_net ), 
        .I2C0_SCL_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/I2C0_SCL_F2H_SCP_net ), 
        .I2C0_SDA_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/I2C0_SDA_F2H_SCP_net ), 
        .I2C1_BCLK(\SF2Project_MSS_0/MSS_ADLIB_INST/I2C1_BCLK_net ), 
        .I2C1_SCL_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/I2C1_SCL_F2H_SCP_net ), 
        .I2C1_SDA_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/I2C1_SDA_F2H_SCP_net ), .MDIF(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDIF_net ), .MGPIO0A_F2H_GPIN(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO0A_F2H_GPIN_net ), 
        .MGPIO10A_F2H_GPIN(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO10A_F2H_GPIN_net ), 
        .MGPIO11A_F2H_GPIN(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO11A_F2H_GPIN_net ), 
        .MGPIO11B_F2H_GPIN(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO11B_F2H_GPIN_net ), 
        .MGPIO12A_F2H_GPIN(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO12A_F2H_GPIN_net ), 
        .MGPIO13A_F2H_GPIN(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO13A_F2H_GPIN_net ), 
        .MGPIO14A_F2H_GPIN(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO14A_F2H_GPIN_net ), 
        .MGPIO15A_F2H_GPIN(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO15A_F2H_GPIN_net ), 
        .MGPIO16A_F2H_GPIN(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO16A_F2H_GPIN_net ), 
        .MGPIO17B_F2H_GPIN(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO17B_F2H_GPIN_net ), 
        .MGPIO18B_F2H_GPIN(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO18B_F2H_GPIN_net ), 
        .MGPIO19B_F2H_GPIN(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO19B_F2H_GPIN_net ), 
        .MGPIO1A_F2H_GPIN(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO1A_F2H_GPIN_net ), 
        .MGPIO20B_F2H_GPIN(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO20B_F2H_GPIN_net ), 
        .MGPIO21B_F2H_GPIN(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO21B_F2H_GPIN_net ), 
        .MGPIO22B_F2H_GPIN(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO22B_F2H_GPIN_net ), 
        .MGPIO24B_F2H_GPIN(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO24B_F2H_GPIN_net ), 
        .MGPIO25B_F2H_GPIN(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO25B_F2H_GPIN_net ), 
        .MGPIO26B_F2H_GPIN(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO26B_F2H_GPIN_net ), 
        .MGPIO27B_F2H_GPIN(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO27B_F2H_GPIN_net ), 
        .MGPIO28B_F2H_GPIN(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO28B_F2H_GPIN_net ), 
        .MGPIO29B_F2H_GPIN(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO29B_F2H_GPIN_net ), 
        .MGPIO2A_F2H_GPIN(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO2A_F2H_GPIN_net ), 
        .MGPIO30B_F2H_GPIN(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO30B_F2H_GPIN_net ), 
        .MGPIO31B_F2H_GPIN(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO31B_F2H_GPIN_net ), 
        .MGPIO3A_F2H_GPIN(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO3A_F2H_GPIN_net ), 
        .MGPIO4A_F2H_GPIN(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO4A_F2H_GPIN_net ), 
        .MGPIO5A_F2H_GPIN(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO5A_F2H_GPIN_net ), 
        .MGPIO6A_F2H_GPIN(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO6A_F2H_GPIN_net ), 
        .MGPIO7A_F2H_GPIN(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO7A_F2H_GPIN_net ), 
        .MGPIO8A_F2H_GPIN(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO8A_F2H_GPIN_net ), 
        .MGPIO9A_F2H_GPIN(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO9A_F2H_GPIN_net ), 
        .MMUART0_CTS_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART0_CTS_F2H_SCP_net ), 
        .MMUART0_DCD_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART0_DCD_F2H_SCP_net ), 
        .MMUART0_DSR_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART0_DSR_F2H_SCP_net ), 
        .MMUART0_DTR_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART0_DTR_F2H_SCP_net ), 
        .MMUART0_RI_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART0_RI_F2H_SCP_net ), 
        .MMUART0_RTS_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART0_RTS_F2H_SCP_net ), 
        .MMUART0_RXD_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART0_RXD_F2H_SCP_net ), 
        .MMUART0_SCK_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART0_SCK_F2H_SCP_net ), 
        .MMUART0_TXD_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART0_TXD_F2H_SCP_net ), 
        .MMUART1_CTS_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART1_CTS_F2H_SCP_net ), 
        .MMUART1_DCD_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART1_DCD_F2H_SCP_net ), 
        .MMUART1_DSR_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART1_DSR_F2H_SCP_net ), 
        .MMUART1_RI_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART1_RI_F2H_SCP_net ), 
        .MMUART1_RTS_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART1_RTS_F2H_SCP_net ), 
        .MMUART1_RXD_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART1_RXD_F2H_SCP_net ), 
        .MMUART1_SCK_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART1_SCK_F2H_SCP_net ), 
        .MMUART1_TXD_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART1_TXD_F2H_SCP_net ), 
        .PER2_FABRIC_PRDATA({
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[31] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[30] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[29] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[28] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[27] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[26] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[25] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[24] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[23] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[22] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[21] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[20] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[19] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[18] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[17] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[16] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[15] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[14] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[13] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[12] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[11] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[10] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[9] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[8] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[7] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[6] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[5] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[4] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[0] }), 
        .PER2_FABRIC_PREADY(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PREADY_net ), 
        .PER2_FABRIC_PSLVERR(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PSLVERR_net ), 
        .RCGF({\SF2Project_MSS_0/MSS_ADLIB_INST/RCGF_net[9] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RCGF_net[8] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RCGF_net[7] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RCGF_net[6] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RCGF_net[5] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RCGF_net[4] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RCGF_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RCGF_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RCGF_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RCGF_net[0] }), .RX_CLKPF(
        \SF2Project_MSS_0/MSS_ADLIB_INST/RX_CLKPF_net ), .RX_DVF(
        \SF2Project_MSS_0/MSS_ADLIB_INST/RX_DVF_net ), .RX_ERRF(
        \SF2Project_MSS_0/MSS_ADLIB_INST/RX_ERRF_net ), .RX_EV(
        \SF2Project_MSS_0/MSS_ADLIB_INST/RX_EV_net ), .RXDF({
        \SF2Project_MSS_0/MSS_ADLIB_INST/RXDF_net[7] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RXDF_net[6] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RXDF_net[5] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RXDF_net[4] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RXDF_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RXDF_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RXDF_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/RXDF_net[0] }), .SLEEPHOLDREQ(
        \SF2Project_MSS_0/MSS_ADLIB_INST/SLEEPHOLDREQ_net ), 
        .SMBALERT_NI0(
        \SF2Project_MSS_0/MSS_ADLIB_INST/SMBALERT_NI0_net ), 
        .SMBALERT_NI1(
        \SF2Project_MSS_0/MSS_ADLIB_INST/SMBALERT_NI1_net ), 
        .SMBSUS_NI0(\SF2Project_MSS_0/MSS_ADLIB_INST/SMBSUS_NI0_net ), 
        .SMBSUS_NI1(\SF2Project_MSS_0/MSS_ADLIB_INST/SMBSUS_NI1_net ), 
        .SPI0_CLK_IN(\SF2Project_MSS_0/MSS_ADLIB_INST/SPI0_CLK_IN_net )
        , .SPI0_SDI_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI0_SDI_F2H_SCP_net ), 
        .SPI0_SDO_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI0_SDO_F2H_SCP_net ), 
        .SPI0_SS0_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI0_SS0_F2H_SCP_net ), 
        .SPI0_SS1_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI0_SS1_F2H_SCP_net ), 
        .SPI0_SS2_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI0_SS2_F2H_SCP_net ), 
        .SPI0_SS3_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI0_SS3_F2H_SCP_net ), 
        .SPI1_CLK_IN(\SF2Project_MSS_0/MSS_ADLIB_INST/SPI1_CLK_IN_net )
        , .SPI1_SDI_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI1_SDI_F2H_SCP_net ), 
        .SPI1_SDO_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI1_SDO_F2H_SCP_net ), 
        .SPI1_SS0_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI1_SS0_F2H_SCP_net ), 
        .SPI1_SS1_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI1_SS1_F2H_SCP_net ), 
        .SPI1_SS2_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI1_SS2_F2H_SCP_net ), 
        .SPI1_SS3_F2H_SCP(
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI1_SS3_F2H_SCP_net ), 
        .TX_CLKPF(\SF2Project_MSS_0/MSS_ADLIB_INST/TX_CLKPF_net ), 
        .USER_MSS_GPIO_RESET_N(
        \SF2Project_MSS_0/MSS_ADLIB_INST/USER_MSS_GPIO_RESET_N_net ), 
        .USER_MSS_RESET_N(
        \SF2Project_MSS_0/MSS_ADLIB_INST/USER_MSS_RESET_N_net ), 
        .XCLK_FAB(\SF2Project_MSS_0/MSS_ADLIB_INST/XCLK_FAB_net ), 
        .CLK_BASE(\SF2Project_MSS_0/MSS_ADLIB_INST/CLK_BASE_net ), 
        .CLK_MDDR_APB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/CLK_MDDR_APB_net ), 
        .F_ARADDR_HADDR1({
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[31] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[30] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[29] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[28] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[27] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[26] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[25] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[24] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[23] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[22] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[21] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[20] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[19] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[18] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[17] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[16] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[15] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[14] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[13] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[12] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[11] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[10] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[9] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[8] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[7] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[6] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[5] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[4] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[0] }), 
        .F_ARBURST_HTRANS1({
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARBURST_HTRANS1_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARBURST_HTRANS1_net[0] }), 
        .F_ARID_HSEL1({
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[0] }), 
        .F_ARLEN_HBURST1({
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[0] }), 
        .F_ARLOCK_HMASTLOCK1({
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARLOCK_HMASTLOCK1_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARLOCK_HMASTLOCK1_net[0] }), 
        .F_ARSIZE_HSIZE1({
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARSIZE_HSIZE1_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARSIZE_HSIZE1_net[0] }), 
        .F_ARVALID_HWRITE1(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARVALID_HWRITE1_net ), 
        .F_AWADDR_HADDR0({
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[31] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[30] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[29] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[28] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[27] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[26] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[25] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[24] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[23] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[22] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[21] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[20] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[19] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[18] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[17] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[16] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[15] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[14] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[13] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[12] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[11] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[10] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[9] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[8] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[7] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[6] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[5] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[4] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[0] }), 
        .F_AWBURST_HTRANS0({
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWBURST_HTRANS0_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWBURST_HTRANS0_net[0] }), 
        .F_AWID_HSEL0({
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[0] }), 
        .F_AWLEN_HBURST0({
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[0] }), 
        .F_AWLOCK_HMASTLOCK0({
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWLOCK_HMASTLOCK0_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWLOCK_HMASTLOCK0_net[0] }), 
        .F_AWSIZE_HSIZE0({
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWSIZE_HSIZE0_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWSIZE_HSIZE0_net[0] }), 
        .F_AWVALID_HWRITE0(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWVALID_HWRITE0_net ), 
        .F_BREADY(\SF2Project_MSS_0/MSS_ADLIB_INST/F_BREADY_net ), 
        .F_RMW_AXI(\SF2Project_MSS_0/MSS_ADLIB_INST/F_RMW_AXI_net ), 
        .F_RREADY(\SF2Project_MSS_0/MSS_ADLIB_INST/F_RREADY_net ), 
        .F_WDATA_HWDATA01({
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[63] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[62] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[61] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[60] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[59] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[58] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[57] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[56] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[55] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[54] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[53] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[52] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[51] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[50] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[49] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[48] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[47] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[46] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[45] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[44] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[43] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[42] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[41] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[40] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[39] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[38] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[37] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[36] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[35] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[34] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[33] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[32] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[31] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[30] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[29] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[28] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[27] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[26] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[25] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[24] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[23] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[22] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[21] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[20] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[19] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[18] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[17] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[16] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[15] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[14] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[13] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[12] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[11] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[10] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[9] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[8] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[7] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[6] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[5] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[4] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[0] }), 
        .F_WID_HREADY01({
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[0] }), 
        .F_WLAST(\SF2Project_MSS_0/MSS_ADLIB_INST/F_WLAST_net ), 
        .F_WSTRB({\SF2Project_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[7] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[6] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[5] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[4] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[0] }), .F_WVALID(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WVALID_net ), 
        .FPGA_MDDR_ARESET_N(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FPGA_MDDR_ARESET_N_net ), 
        .MDDR_FABRIC_PADDR({
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[10] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[9] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[8] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[7] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[6] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[5] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[4] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[2] }), 
        .MDDR_FABRIC_PENABLE(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PENABLE_net ), 
        .MDDR_FABRIC_PSEL(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PSEL_net ), 
        .MDDR_FABRIC_PWDATA({
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[15] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[14] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[13] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[12] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[11] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[10] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[9] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[8] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[7] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[6] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[5] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[4] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[3] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[2] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[1] , 
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[0] }), 
        .MDDR_FABRIC_PWRITE(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWRITE_net ), 
        .PRESET_N(\SF2Project_MSS_0/MSS_ADLIB_INST/PRESET_N_net ), 
        .CAN_RXBUS_USBA_DATA1_MGPIO3A_IN(GND), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN(GND), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_IN(GND), .DM_IN({GND, 
        \SF2Project_MSS_0/MDDR_DM_RDQS_1_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DM_RDQS_0_PAD_Y }), .DRAM_DQ_IN({GND, 
        GND, \SF2Project_MSS_0/MDDR_DQ_15_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DQ_14_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DQ_13_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DQ_12_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DQ_11_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DQ_10_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DQ_9_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DQ_8_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DQ_7_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DQ_6_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DQ_5_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DQ_4_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DQ_3_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DQ_2_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DQ_1_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DQ_0_PAD_Y }), .DRAM_DQS_IN({GND, 
        \SF2Project_MSS_0/MDDR_DQS_1_PAD_Y , 
        \SF2Project_MSS_0/MDDR_DQS_0_PAD_Y }), .DRAM_FIFO_WE_IN({GND, 
        \SF2Project_MSS_0/MDDR_DQS_TMATCH_0_IN_PAD_Y }), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_IN(
        \SF2Project_MSS_0/I2C_0_SCL_PAD_Y ), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_IN(
        \SF2Project_MSS_0/I2C_0_SDA_PAD_Y ), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_IN(
        \SF2Project_MSS_0/I2C_1_SCL_PAD_Y ), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_IN(
        \SF2Project_MSS_0/I2C_1_SDA_PAD_Y ), 
        .MMUART0_CTS_USBC_DATA7_MGPIO19B_IN(GND), 
        .MMUART0_DCD_MGPIO22B_IN(GND), .MMUART0_DSR_MGPIO20B_IN(GND), 
        .MMUART0_DTR_USBC_DATA6_MGPIO18B_IN(GND), 
        .MMUART0_RI_MGPIO21B_IN(GND), 
        .MMUART0_RTS_USBC_DATA5_MGPIO17B_IN(GND), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_IN(
        \SF2Project_MSS_0/MMUART_0_RXD_PAD_Y ), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_IN(GND), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_IN(GND), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_IN(
        \SF2Project_MSS_0/MMUART_1_RXD_PAD_Y ), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_IN(GND), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_IN(GND), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN(
        \SF2Project_MSS_0/USB_ULPI_XCLK_PAD_Y ), 
        .RGMII_MDC_RMII_MDC_IN(GND), 
        .RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN(
        \SF2Project_MSS_0/USB_ULPI_DATA_7_PAD_Y ), .RGMII_RX_CLK_IN(
        GND), .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN(
        \SF2Project_MSS_0/USB_ULPI_DATA_2_PAD_Y ), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN(
        \SF2Project_MSS_0/USB_ULPI_DATA_0_PAD_Y ), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN(
        \SF2Project_MSS_0/USB_ULPI_DATA_1_PAD_Y ), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN(
        \SF2Project_MSS_0/USB_ULPI_DATA_3_PAD_Y ), 
        .RGMII_RXD3_USBB_DATA4_IN(
        \SF2Project_MSS_0/USB_ULPI_DATA_4_PAD_Y ), .RGMII_TX_CLK_IN(
        GND), .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN(
        \SF2Project_MSS_0/USB_ULPI_NXT_PAD_Y ), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_IN(
        \SF2Project_MSS_0/USB_ULPI_DIR_PAD_Y ), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_IN(GND), 
        .RGMII_TXD2_USBB_DATA5_IN(
        \SF2Project_MSS_0/USB_ULPI_DATA_5_PAD_Y ), 
        .RGMII_TXD3_USBB_DATA6_IN(
        \SF2Project_MSS_0/USB_ULPI_DATA_6_PAD_Y ), 
        .SPI0_SCK_USBA_XCLK_IN(\SF2Project_MSS_0/SPI_0_CLK_PAD_Y ), 
        .SPI0_SDI_USBA_DIR_MGPIO5A_IN(
        \SF2Project_MSS_0/SPI_0_DI_PAD_Y ), 
        .SPI0_SDO_USBA_STP_MGPIO6A_IN(GND), 
        .SPI0_SS0_USBA_NXT_MGPIO7A_IN(
        \SF2Project_MSS_0/SPI_0_SS0_PAD_Y ), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_IN(GND), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_IN(GND), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_IN(GND), .SPI1_SCK_IN(
        \SF2Project_MSS_0/SPI_1_CLK_PAD_Y ), .SPI1_SDI_MGPIO11A_IN(
        \SF2Project_MSS_0/SPI_1_DI_PAD_Y ), .SPI1_SDO_MGPIO12A_IN(GND), 
        .SPI1_SS0_MGPIO13A_IN(\SF2Project_MSS_0/SPI_1_SS0_PAD_Y ), 
        .SPI1_SS1_MGPIO14A_IN(GND), .SPI1_SS2_MGPIO15A_IN(GND), 
        .SPI1_SS3_MGPIO16A_IN(GND), .SPI1_SS4_MGPIO17A_IN(GND), 
        .SPI1_SS5_MGPIO18A_IN(GND), .SPI1_SS6_MGPIO23A_IN(GND), 
        .SPI1_SS7_MGPIO24A_IN(GND), .USBC_XCLK_IN(GND), 
        .CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT(), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT(), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT(), .DRAM_ADDR({
        \SF2Project_MSS_0/DRAM_ADDR_net_0[15] , 
        \SF2Project_MSS_0/DRAM_ADDR_net_0[14] , 
        \SF2Project_MSS_0/DRAM_ADDR_net_0[13] , 
        \SF2Project_MSS_0/DRAM_ADDR_net_0[12] , 
        \SF2Project_MSS_0/DRAM_ADDR_net_0[11] , 
        \SF2Project_MSS_0/DRAM_ADDR_net_0[10] , 
        \SF2Project_MSS_0/DRAM_ADDR_net_0[9] , 
        \SF2Project_MSS_0/DRAM_ADDR_net_0[8] , 
        \SF2Project_MSS_0/DRAM_ADDR_net_0[7] , 
        \SF2Project_MSS_0/DRAM_ADDR_net_0[6] , 
        \SF2Project_MSS_0/DRAM_ADDR_net_0[5] , 
        \SF2Project_MSS_0/DRAM_ADDR_net_0[4] , 
        \SF2Project_MSS_0/DRAM_ADDR_net_0[3] , 
        \SF2Project_MSS_0/DRAM_ADDR_net_0[2] , 
        \SF2Project_MSS_0/DRAM_ADDR_net_0[1] , 
        \SF2Project_MSS_0/DRAM_ADDR_net_0[0] }), .DRAM_BA({
        \SF2Project_MSS_0/DRAM_BA_net_0[2] , 
        \SF2Project_MSS_0/DRAM_BA_net_0[1] , 
        \SF2Project_MSS_0/DRAM_BA_net_0[0] }), .DRAM_CASN(
        \SF2Project_MSS_0/MSS_ADLIB_INST_DRAM_CASN ), .DRAM_CKE(
        \SF2Project_MSS_0/MSS_ADLIB_INST_DRAM_CKE ), .DRAM_CLK(
        \SF2Project_MSS_0/MSS_ADLIB_INST_DRAM_CLK ), .DRAM_CSN(
        \SF2Project_MSS_0/MSS_ADLIB_INST_DRAM_CSN ), .DRAM_DM_RDQS_OUT({
        nc302, \SF2Project_MSS_0/DRAM_DM_RDQS_OUT_net_0[1] , 
        \SF2Project_MSS_0/DRAM_DM_RDQS_OUT_net_0[0] }), .DRAM_DQ_OUT({
        nc303, nc304, \SF2Project_MSS_0/DRAM_DQ_OUT_net_0[15] , 
        \SF2Project_MSS_0/DRAM_DQ_OUT_net_0[14] , 
        \SF2Project_MSS_0/DRAM_DQ_OUT_net_0[13] , 
        \SF2Project_MSS_0/DRAM_DQ_OUT_net_0[12] , 
        \SF2Project_MSS_0/DRAM_DQ_OUT_net_0[11] , 
        \SF2Project_MSS_0/DRAM_DQ_OUT_net_0[10] , 
        \SF2Project_MSS_0/DRAM_DQ_OUT_net_0[9] , 
        \SF2Project_MSS_0/DRAM_DQ_OUT_net_0[8] , 
        \SF2Project_MSS_0/DRAM_DQ_OUT_net_0[7] , 
        \SF2Project_MSS_0/DRAM_DQ_OUT_net_0[6] , 
        \SF2Project_MSS_0/DRAM_DQ_OUT_net_0[5] , 
        \SF2Project_MSS_0/DRAM_DQ_OUT_net_0[4] , 
        \SF2Project_MSS_0/DRAM_DQ_OUT_net_0[3] , 
        \SF2Project_MSS_0/DRAM_DQ_OUT_net_0[2] , 
        \SF2Project_MSS_0/DRAM_DQ_OUT_net_0[1] , 
        \SF2Project_MSS_0/DRAM_DQ_OUT_net_0[0] }), .DRAM_DQS_OUT({
        nc305, \SF2Project_MSS_0/DRAM_DQS_OUT_net_0[1] , 
        \SF2Project_MSS_0/DRAM_DQS_OUT_net_0[0] }), .DRAM_FIFO_WE_OUT({
        nc306, \SF2Project_MSS_0/DRAM_FIFO_WE_OUT_net_0[0] }), 
        .DRAM_ODT(\SF2Project_MSS_0/MSS_ADLIB_INST_DRAM_ODT ), 
        .DRAM_RASN(\SF2Project_MSS_0/MSS_ADLIB_INST_DRAM_RASN ), 
        .DRAM_RSTN(\SF2Project_MSS_0/MSS_ADLIB_INST_DRAM_RSTN ), 
        .DRAM_WEN(\SF2Project_MSS_0/MSS_ADLIB_INST_DRAM_WEN ), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_OUT(
        \SF2Project_MSS_0/MSS_ADLIB_INST_I2C0_SCL_USBC_DATA1_MGPIO31B_OUT )
        , .I2C0_SDA_USBC_DATA0_MGPIO30B_OUT(
        \SF2Project_MSS_0/MSS_ADLIB_INST_I2C0_SDA_USBC_DATA0_MGPIO30B_OUT )
        , .I2C1_SCL_USBA_DATA4_MGPIO1A_OUT(
        \SF2Project_MSS_0/MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OUT )
        , .I2C1_SDA_USBA_DATA3_MGPIO0A_OUT(
        \SF2Project_MSS_0/MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OUT )
        , .MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT(), 
        .MMUART0_DCD_MGPIO22B_OUT(), .MMUART0_DSR_MGPIO20B_OUT(), 
        .MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT(), 
        .MMUART0_RI_MGPIO21B_OUT(), 
        .MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT(), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_OUT(), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_OUT(), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_OUT(
        \SF2Project_MSS_0/MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OUT )
        , .MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT(), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT(), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT(
        \SF2Project_MSS_0/MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT )
        , .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT(), 
        .RGMII_MDC_RMII_MDC_OUT(), 
        .RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT(
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT )
        , .RGMII_RX_CLK_OUT(), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT(
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT )
        , .RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT(
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT )
        , .RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT(
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT )
        , .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT(
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT )
        , .RGMII_RXD3_USBB_DATA4_OUT(
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_RXD3_USBB_DATA4_OUT ), 
        .RGMII_TX_CLK_OUT(), .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT(), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT(), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_OUT(
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_TXD1_RMII_TXD1_USBB_STP_OUT )
        , .RGMII_TXD2_USBB_DATA5_OUT(
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_TXD2_USBB_DATA5_OUT ), 
        .RGMII_TXD3_USBB_DATA6_OUT(
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_TXD3_USBB_DATA6_OUT ), 
        .SPI0_SCK_USBA_XCLK_OUT(
        \SF2Project_MSS_0/MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OUT ), 
        .SPI0_SDI_USBA_DIR_MGPIO5A_OUT(), 
        .SPI0_SDO_USBA_STP_MGPIO6A_OUT(
        \SF2Project_MSS_0/MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OUT )
        , .SPI0_SS0_USBA_NXT_MGPIO7A_OUT(
        \SF2Project_MSS_0/MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OUT )
        , .SPI0_SS1_USBA_DATA5_MGPIO8A_OUT(), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_OUT(), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_OUT(), .SPI1_SCK_OUT(
        \SF2Project_MSS_0/MSS_ADLIB_INST_SPI1_SCK_OUT ), 
        .SPI1_SDI_MGPIO11A_OUT(), .SPI1_SDO_MGPIO12A_OUT(
        \SF2Project_MSS_0/MSS_ADLIB_INST_SPI1_SDO_MGPIO12A_OUT ), 
        .SPI1_SS0_MGPIO13A_OUT(
        \SF2Project_MSS_0/MSS_ADLIB_INST_SPI1_SS0_MGPIO13A_OUT ), 
        .SPI1_SS1_MGPIO14A_OUT(), .SPI1_SS2_MGPIO15A_OUT(), 
        .SPI1_SS3_MGPIO16A_OUT(), .SPI1_SS4_MGPIO17A_OUT(), 
        .SPI1_SS5_MGPIO18A_OUT(), .SPI1_SS6_MGPIO23A_OUT(), 
        .SPI1_SS7_MGPIO24A_OUT(), .USBC_XCLK_OUT(), 
        .CAN_RXBUS_USBA_DATA1_MGPIO3A_OE(), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE(), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_OE(), .DM_OE({nc307, 
        \SF2Project_MSS_0/DM_OE_net_0[1] , 
        \SF2Project_MSS_0/DM_OE_net_0[0] }), .DRAM_DQ_OE({nc308, nc309, 
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[15] , 
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[14] , 
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[13] , 
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[12] , 
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[11] , 
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[10] , 
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[9] , 
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[8] , 
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[7] , 
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[6] , 
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[5] , 
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[4] , 
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[3] , 
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[2] , 
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[1] , 
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[0] }), .DRAM_DQS_OE({nc310, 
        \SF2Project_MSS_0/DRAM_DQS_OE_net_0[1] , 
        \SF2Project_MSS_0/DRAM_DQS_OE_net_0[0] }), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_OE(
        \SF2Project_MSS_0/MSS_ADLIB_INST_I2C0_SCL_USBC_DATA1_MGPIO31B_OE )
        , .I2C0_SDA_USBC_DATA0_MGPIO30B_OE(
        \SF2Project_MSS_0/MSS_ADLIB_INST_I2C0_SDA_USBC_DATA0_MGPIO30B_OE )
        , .I2C1_SCL_USBA_DATA4_MGPIO1A_OE(
        \SF2Project_MSS_0/MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OE )
        , .I2C1_SDA_USBA_DATA3_MGPIO0A_OE(
        \SF2Project_MSS_0/MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OE )
        , .MMUART0_CTS_USBC_DATA7_MGPIO19B_OE(), 
        .MMUART0_DCD_MGPIO22B_OE(), .MMUART0_DSR_MGPIO20B_OE(), 
        .MMUART0_DTR_USBC_DATA6_MGPIO18B_OE(), .MMUART0_RI_MGPIO21B_OE(
        ), .MMUART0_RTS_USBC_DATA5_MGPIO17B_OE(), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_OE(), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_OE(), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_OE(
        \SF2Project_MSS_0/MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OE )
        , .MMUART1_RXD_USBC_DATA3_MGPIO26B_OE(), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_OE(), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_OE(
        \SF2Project_MSS_0/MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OE )
        , .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE(), 
        .RGMII_MDC_RMII_MDC_OE(), .RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE(
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE )
        , .RGMII_RX_CLK_OE(), .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE(
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE )
        , .RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE(
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE )
        , .RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE(
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE )
        , .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE(
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE )
        , .RGMII_RXD3_USBB_DATA4_OE(
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_RXD3_USBB_DATA4_OE ), 
        .RGMII_TX_CLK_OE(), .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE(), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_OE(), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_OE(
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_TXD1_RMII_TXD1_USBB_STP_OE )
        , .RGMII_TXD2_USBB_DATA5_OE(
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_TXD2_USBB_DATA5_OE ), 
        .RGMII_TXD3_USBB_DATA6_OE(
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_TXD3_USBB_DATA6_OE ), 
        .SPI0_SCK_USBA_XCLK_OE(
        \SF2Project_MSS_0/MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OE ), 
        .SPI0_SDI_USBA_DIR_MGPIO5A_OE(), .SPI0_SDO_USBA_STP_MGPIO6A_OE(
        \SF2Project_MSS_0/MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OE )
        , .SPI0_SS0_USBA_NXT_MGPIO7A_OE(
        \SF2Project_MSS_0/MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OE )
        , .SPI0_SS1_USBA_DATA5_MGPIO8A_OE(), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_OE(), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_OE(), .SPI1_SCK_OE(
        \SF2Project_MSS_0/MSS_ADLIB_INST_SPI1_SCK_OE ), 
        .SPI1_SDI_MGPIO11A_OE(), .SPI1_SDO_MGPIO12A_OE(
        \SF2Project_MSS_0/MSS_ADLIB_INST_SPI1_SDO_MGPIO12A_OE ), 
        .SPI1_SS0_MGPIO13A_OE(
        \SF2Project_MSS_0/MSS_ADLIB_INST_SPI1_SS0_MGPIO13A_OE ), 
        .SPI1_SS1_MGPIO14A_OE(), .SPI1_SS2_MGPIO15A_OE(), 
        .SPI1_SS3_MGPIO16A_OE(), .SPI1_SS4_MGPIO17A_OE(), 
        .SPI1_SS5_MGPIO18A_OE(), .SPI1_SS6_MGPIO23A_OE(), 
        .SPI1_SS7_MGPIO24A_OE(), .USBC_XCLK_OE());
    sdf_IOPAD_BI \SF2Project_MSS_0/MDDR_DQ_2_PAD/U_IOPAD  (.PAD(
        MDDR_DQ[2]), .D(\SF2Project_MSS_0/DRAM_DQ_OUT_net_0[2] ), .E(
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[2] ), .Y(
        \SF2Project_MSS_0/MDDR_DQ_2_PAD_Y ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_87  (.A(
        VCC), .B(\MAC_MII_RXD[3] ), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[28] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/RXDF_net[3] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_169  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART1_DSR_F2H_SCP_net ), 
        .IPB(), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_36  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[19] ), .IPB(), 
        .IPC());
    IOBI_IB_OB_EB \SF2Project_MSS_0/I2C_1_SDA_PAD/U_IOBI  (.D(VCC), .E(
        VCC), .YIN(\SF2Project_MSS_0/I2C_1_SDA_PAD/YIN ), .DOUT(), 
        .EOUT(), .Y());
    IOTRI_OB_EB \SF2Project_MSS_0/USB_ULPI_STP_PAD/U_IOOUT  (.D(VCC), 
        .E(VCC), .DOUT(), .EOUT());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_253  (
        .A(VCC), .B(VCC), .C(GND), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[1] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[13] )
        , .IPC(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARSIZE_HSIZE1_net[1] ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_160  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO11A_F2H_GPIN_net ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO14A_F2H_GPIN_net ), .IPC(
        ));
    IOINFF_BYPASS \SF2Project_MSS_0/MDDR_DQ_9_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/MDDR_DQ_9_PAD_Y ), .Y(
        \SF2Project_MSS_0/MDDR_DQ_9_PAD/YIN ));
    IOIN_IB \SF2Project_MSS_0/MDDR_DQS_1_PAD/U_IOP  (.YIN(
        \SF2Project_MSS_0/MDDR_DQS_1_PAD/YIN ), .E(GND), .Y());
    IOTRI_OB_EB \SF2Project_MSS_0/SPI_0_DO_PAD/U_IOOUT  (.D(VCC), .E(
        VCC), .DOUT(), .EOUT());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_213  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[31] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[1] ), 
        .IPC());
    sdf_IOPAD_BI \SF2Project_MSS_0/I2C_0_SDA_PAD/U_IOPAD  (.PAD(
        I2C_0_SDA), .D(
        \SF2Project_MSS_0/MSS_ADLIB_INST_I2C0_SDA_USBC_DATA0_MGPIO30B_OUT )
        , .E(
        \SF2Project_MSS_0/MSS_ADLIB_INST_I2C0_SDA_USBC_DATA0_MGPIO30B_OE )
        , .Y(\SF2Project_MSS_0/I2C_0_SDA_PAD_Y ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_251  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[63] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[3] ), 
        .IPC());
    IOINFF_BYPASS \SF2Project_MSS_0/MDDR_DQ_13_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/MDDR_DQ_13_PAD_Y ), .Y(
        \SF2Project_MSS_0/MDDR_DQ_13_PAD/YIN ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_211  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[29] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWLOCK_HMASTLOCK0_net[1] ), 
        .IPC());
    sdf_IOPAD_TRI \SF2Project_MSS_0/MDDR_BA_0_PAD/U_IOPAD  (.PAD(
        MDDR_BA[0]), .D(\SF2Project_MSS_0/DRAM_BA_net_0[0] ), .E(
        \SF2Project_MSS_0/MDDR_BA_0_PAD/EOUT ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_86  (.A(
        VCC), .B(\MAC_MII_RXD[2] ), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[27] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/RXDF_net[2] ), .IPC());
    CFG1 #( .INIT(2'h2) )  BLOCK_INTERFACE_I_MAC_MII_RX_DV (.A(
        MAC_MII_RX_DV), .Y(MAC_MII_RX_DV_net_1));
    IOINFF_BYPASS \SF2Project_MSS_0/USB_ULPI_DATA_3_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/USB_ULPI_DATA_3_PAD_Y ), .Y(
        \SF2Project_MSS_0/USB_ULPI_DATA_3_PAD/YIN ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_257  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[5] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[17] )
        , .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_217  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[1] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[13] ), 
        .IPC(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[25] ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_229  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[27] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[39] ), 
        .IPC(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[51] ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_239  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[37] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[49] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_19  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[24] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[31] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_12  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[17] ), .IPB(), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_4  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[2] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[9] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_206  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[24] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[2] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_13  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[18] ), .IPB(), 
        .IPC());
    sdf_IOPAD_TRI \SF2Project_MSS_0/MDDR_ADDR_8_PAD/U_IOPAD  (.PAD(
        MDDR_ADDR[8]), .D(\SF2Project_MSS_0/DRAM_ADDR_net_0[8] ), .E(
        \SF2Project_MSS_0/MDDR_ADDR_8_PAD/EOUT ));
    IOINFF_BYPASS \SF2Project_MSS_0/I2C_1_SCL_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/I2C_1_SCL_PAD_Y ), .Y(
        \SF2Project_MSS_0/I2C_1_SCL_PAD/YIN ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_148  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO1A_F2H_GPIN_net ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/CAN_TX_EBL_F2H_SCP_net ), 
        .IPC());
    CFG1 #( .INIT(2'h2) )  BLOCK_INTERFACE_I_MAC_MII_RX_CLK (.A(
        MAC_MII_RX_CLK), .Y(MAC_MII_RX_CLK_net_1));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_273  (
        .A(GND), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[1] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PSEL_net ), 
        .IPC());
    IOTRI_OB_EB \SF2Project_MSS_0/MDDR_ADDR_8_PAD/U_IOOUT  (.D(VCC), 
        .E(VCC), .DOUT(), .EOUT(
        \SF2Project_MSS_0/MDDR_ADDR_8_PAD/EOUT ));
    IOBI_IB_OB_EB \SF2Project_MSS_0/USB_ULPI_DATA_2_PAD/U_IOBI  (.D(
        VCC), .E(VCC), .YIN(\SF2Project_MSS_0/USB_ULPI_DATA_2_PAD/YIN )
        , .DOUT(), .EOUT(), .Y());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_271  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[31] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/FPGA_MDDR_ARESET_N_net ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_200  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[4] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[16] )
        , .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_194  (
        .A(GND), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[2] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[10] ), 
        .IPC());
    sdf_IOPADN_TRI \SF2Project_MSS_0/MDDR_CLK_PAD/U_IOPADN  (.PAD_P(
        MDDR_CLK_N), .OIN_P(\SF2Project_MSS_0/MSS_ADLIB_INST_DRAM_CLK )
        , .EIN_P(VCC));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_59  (.A(
        VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[20] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_224  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[8] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[20] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_124  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_IDDIG_net ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[6] ), .IPC()
        );
    sdf_IOPAD_BI \SF2Project_MSS_0/MDDR_DQ_11_PAD/U_IOPAD  (.PAD(
        MDDR_DQ[11]), .D(\SF2Project_MSS_0/DRAM_DQ_OUT_net_0[11] ), .E(
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[11] ), .Y(
        \SF2Project_MSS_0/MDDR_DQ_11_PAD_Y ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_52  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[6] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[13] ), .IPC());
    IOTRI_OB_EB \SF2Project_MSS_0/MDDR_CS_N_PAD/U_IOOUT  (.D(VCC), .E(
        VCC), .DOUT(), .EOUT(\SF2Project_MSS_0/MDDR_CS_N_PAD/EOUT ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_255  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[3] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[15] )
        , .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_234  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[32] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[44] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_134  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/I2C0_BCLK_net ), .IPB(), .IPC(
        ));
    sdf_IOPAD_IN \SF2Project_MSS_0/USB_ULPI_XCLK_PAD/U_IOPAD  (.PAD(
        USB_ULPI_XCLK), .Y(\SF2Project_MSS_0/USB_ULPI_XCLK_PAD_Y ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_53  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[7] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[14] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_215  (
        .A(GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWSIZE_HSIZE0_net[1] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[3] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_277  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[1] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[4] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_199  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[3] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[15] )
        , .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_188  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO30B_F2H_GPIN_net ), .IPB(
        ), .IPC());
    sdf_IOPAD_BI \SF2Project_MSS_0/SPI_0_SS0_PAD/U_IOPAD  (.PAD(
        SPI_0_SS0), .D(
        \SF2Project_MSS_0/MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OUT )
        , .E(
        \SF2Project_MSS_0/MSS_ADLIB_INST_SPI0_SS0_USBA_NXT_MGPIO7A_OE )
        , .Y(\SF2Project_MSS_0/SPI_0_SS0_PAD_Y ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_39  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[22] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[29] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_129  (
        .A(GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[4] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[11] ), .IPC(
        ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_32  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[8] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[15] ), .IPC());
    IOBI_IB_OB_EB \SF2Project_MSS_0/USB_ULPI_DATA_5_PAD/U_IOBI  (.D(
        VCC), .E(VCC), .YIN(\SF2Project_MSS_0/USB_ULPI_DATA_5_PAD/YIN )
        , .DOUT(), .EOUT(), .Y());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_139  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/SMBSUS_NI1_net ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2_DMAREADY_net[1] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_44  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[27] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_READY_net ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_33  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[9] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[16] ), .IPC());
    IOINFF_BYPASS \SF2Project_MSS_0/USB_ULPI_DATA_5_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/USB_ULPI_DATA_5_PAD_Y ), .Y(
        \SF2Project_MSS_0/USB_ULPI_DATA_5_PAD/YIN ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_263  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[11] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[23] )
        , .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_120  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_VBUSVALID_net ), .IPB(), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_261  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[9] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[21] )
        , .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_130  (
        .A(VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[12] ), .IPC(
        ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_0  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_READY_net ), .IPB(), 
        .IPC());
    IOINFF_BYPASS \SF2Project_MSS_0/MDDR_DQ_12_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/MDDR_DQ_12_PAD_Y ), .Y(
        \SF2Project_MSS_0/MDDR_DQ_12_PAD/YIN ));
    sdf_IOPAD_TRI \SF2Project_MSS_0/MDDR_RAS_N_PAD/U_IOPAD  (.PAD(
        MDDR_RAS_N), .D(\SF2Project_MSS_0/MSS_ADLIB_INST_DRAM_RASN ), 
        .E(\SF2Project_MSS_0/MDDR_RAS_N_PAD/EOUT ));
    sdf_IOPAD_BI \SF2Project_MSS_0/MDDR_DQ_3_PAD/U_IOPAD  (.PAD(
        MDDR_DQ[3]), .D(\SF2Project_MSS_0/DRAM_DQ_OUT_net_0[3] ), .E(
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[3] ), .Y(
        \SF2Project_MSS_0/MDDR_DQ_3_PAD_Y ));
    IOINFF_BYPASS \SF2Project_MSS_0/MDDR_DQ_11_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/MDDR_DQ_11_PAD_Y ), .Y(
        \SF2Project_MSS_0/MDDR_DQ_11_PAD/YIN ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_89  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[30] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/RXDF_net[5] ), .IPC());
    sdf_IOPAD_BI \SF2Project_MSS_0/MDDR_DQ_5_PAD/U_IOPAD  (.PAD(
        MDDR_DQ[5]), .D(\SF2Project_MSS_0/DRAM_DQ_OUT_net_0[5] ), .E(
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[5] ), .Y(
        \SF2Project_MSS_0/MDDR_DQ_5_PAD_Y ));
    sdf_IOPAD_BI \SF2Project_MSS_0/USB_ULPI_DATA_2_PAD/U_IOPAD  (.PAD(
        USB_ULPI_DATA[2]), .D(
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT )
        , .E(
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE )
        , .Y(\SF2Project_MSS_0/USB_ULPI_DATA_2_PAD_Y ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_82  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[23] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_70  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[4] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_267  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[27] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARLOCK_HMASTLOCK1_net[1] ), 
        .IPC());
    IOBI_IB_OB_EB \SF2Project_MSS_0/MDDR_DQ_8_PAD/U_IOBI  (.D(VCC), .E(
        VCC), .YIN(\SF2Project_MSS_0/MDDR_DQ_8_PAD/YIN ), .DOUT(), 
        .EOUT(), .Y());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_83  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[24] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_101  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/RCGF_net[1] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/RCGF_net[8] ), .IPC());
    IOBI_IB_OB_EB \SF2Project_MSS_0/USB_ULPI_DATA_3_PAD/U_IOBI  (.D(
        VCC), .E(VCC), .YIN(\SF2Project_MSS_0/USB_ULPI_DATA_3_PAD/YIN )
        , .DOUT(), .EOUT(), .Y());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_48  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[2] ), .IPB(), 
        .IPC());
    sdf_IOPAD_TRI \SF2Project_MSS_0/MDDR_ADDR_12_PAD/U_IOPAD  (.PAD(
        MDDR_ADDR[12]), .D(\SF2Project_MSS_0/DRAM_ADDR_net_0[12] ), .E(
        \SF2Project_MSS_0/MDDR_ADDR_12_PAD/EOUT ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_152  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO3A_F2H_GPIN_net ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI0_SDO_F2H_SCP_net ), .IPC()
        );
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_145  (
        .A(GND), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/SLEEPHOLDREQ_net ), .IPB(), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_112  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[4] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[1] ), .IPC());
    sdf_IOPAD_BI \SF2Project_MSS_0/I2C_0_SCL_PAD/U_IOPAD  (.PAD(
        I2C_0_SCL), .D(
        \SF2Project_MSS_0/MSS_ADLIB_INST_I2C0_SCL_USBC_DATA1_MGPIO31B_OUT )
        , .E(
        \SF2Project_MSS_0/MSS_ADLIB_INST_I2C0_SCL_USBC_DATA1_MGPIO31B_OE )
        , .Y(\SF2Project_MSS_0/I2C_0_SCL_PAD_Y ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_275  (
        .A(GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[3] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/PRESET_N_net ), .IPC());
    IOBI_IB_OB_EB \SF2Project_MSS_0/USB_ULPI_DATA_6_PAD/U_IOBI  (.D(
        VCC), .E(VCC), .YIN(\SF2Project_MSS_0/USB_ULPI_DATA_6_PAD/YIN )
        , .DOUT(), .EOUT(), .Y());
    CFG1 #( .INIT(2'h2) )  BLOCK_INTERFACE_I_MAC_MII_CRS (.A(
        MAC_MII_CRS), .Y(MAC_MII_CRS_net_1));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_106  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_TXREADY_net ), .IPC());
    IOTRI_OB_EB \SF2Project_MSS_0/MDDR_BA_0_PAD/U_IOOUT  (.D(VCC), .E(
        VCC), .DOUT(), .EOUT(\SF2Project_MSS_0/MDDR_BA_0_PAD/EOUT ));
    sdf_IOPAD_IN \SF2Project_MSS_0/SPI_0_DI_PAD/U_IOPAD  (.PAD(
        SPI_0_DI), .Y(\SF2Project_MSS_0/SPI_0_DI_PAD_Y ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_91  (.A(
        MAC_MII_TX_CLK_net_1), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/TX_CLKPF_net ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/RXDF_net[7] ), .IPC());
    IOINFF_BYPASS \SF2Project_MSS_0/MMUART_1_RXD_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/MMUART_1_RXD_PAD_Y ), .Y(
        \SF2Project_MSS_0/MMUART_1_RXD_PAD/YIN ));
    CFG1 #( .INIT(2'h2) )  \BLOCK_INTERFACE_I_MAC_MII_TXD[3]  (.A(
        \MAC_MII_TXD[3] ), .Y(MAC_MII_TXD[3]));
    IOBI_IB_OB_EB \SF2Project_MSS_0/I2C_0_SCL_PAD/U_IOBI  (.D(VCC), .E(
        VCC), .YIN(\SF2Project_MSS_0/I2C_0_SCL_PAD/YIN ), .DOUT(), 
        .EOUT(), .Y());
    CFG1 #( .INIT(2'h2) )  \BLOCK_INTERFACE_I_MAC_MII_TXD[0]  (.A(
        \MAC_MII_TXD[0] ), .Y(MAC_MII_TXD[0]));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_65  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[26] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PSLVERR_net ), 
        .IPC());
    IOTRI_OB_EB \SF2Project_MSS_0/MDDR_ADDR_3_PAD/U_IOOUT  (.D(VCC), 
        .E(VCC), .DOUT(), .EOUT(
        \SF2Project_MSS_0/MDDR_ADDR_3_PAD/EOUT ));
    sdf_IOPAD_TRI \SF2Project_MSS_0/MDDR_ADDR_2_PAD/U_IOPAD  (.PAD(
        MDDR_ADDR[2]), .D(\SF2Project_MSS_0/DRAM_ADDR_net_0[2] ), .E(
        \SF2Project_MSS_0/MDDR_ADDR_2_PAD/EOUT ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_61  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[22] ), .IPB(), 
        .IPC());
    sdf_IOPAD_BI \SF2Project_MSS_0/MDDR_DQ_13_PAD/U_IOPAD  (.PAD(
        MDDR_DQ[13]), .D(\SF2Project_MSS_0/DRAM_DQ_OUT_net_0[13] ), .E(
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[13] ), .Y(
        \SF2Project_MSS_0/MDDR_DQ_13_PAD_Y ));
    IOINFF_BYPASS \SF2Project_MSS_0/MDDR_DQ_0_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/MDDR_DQ_0_PAD_Y ), .Y(
        \SF2Project_MSS_0/MDDR_DQ_0_PAD/YIN ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_185  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART0_RXD_F2H_SCP_net ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/I2C0_SCL_F2H_SCP_net ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_265  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[25] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARBURST_HTRANS1_net[1] ), 
        .IPC(\SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWRITE_net ));
    IOBI_IB_OB_EB \SF2Project_MSS_0/MDDR_DQ_14_PAD/U_IOBI  (.D(VCC), 
        .E(VCC), .YIN(\SF2Project_MSS_0/MDDR_DQ_14_PAD/YIN ), .DOUT(), 
        .EOUT(), .Y());
    sdf_IOPAD_BI \SF2Project_MSS_0/SPI_0_CLK_PAD/U_IOPAD  (.PAD(
        SPI_0_CLK), .D(
        \SF2Project_MSS_0/MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OUT ), .E(
        \SF2Project_MSS_0/MSS_ADLIB_INST_SPI0_SCK_USBA_XCLK_OE ), .Y(
        \SF2Project_MSS_0/SPI_0_CLK_PAD_Y ));
    IOINFF_BYPASS \SF2Project_MSS_0/SPI_0_SS0_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/SPI_0_SS0_PAD_Y ), .Y(
        \SF2Project_MSS_0/SPI_0_SS0_PAD/YIN ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_107  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_RXVALID_net ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_223  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[7] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[19] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_172  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO24B_F2H_GPIN_net ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART0_RTS_F2H_SCP_net ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_103  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/RCGF_net[3] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/XCLK_FAB_net ), .IPC());
    CFG1 #( .INIT(2'h2) )  \BLOCK_INTERFACE_I_MAC_MII_TXD[1]  (.A(
        \MAC_MII_TXD[1] ), .Y(MAC_MII_TXD[1]));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_233  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[31] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[43] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_221  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[5] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[17] ), 
        .IPC());
    IOINFF_BYPASS \SF2Project_MSS_0/MDDR_DM_RDQS_0_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/MDDR_DM_RDQS_0_PAD_Y ), .Y(
        \SF2Project_MSS_0/MDDR_DM_RDQS_0_PAD/YIN ));
    IOTRI_OB_EB \SF2Project_MSS_0/MDDR_BA_2_PAD/U_IOOUT  (.D(VCC), .E(
        VCC), .DOUT(), .EOUT(\SF2Project_MSS_0/MDDR_BA_2_PAD/EOUT ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_231  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[29] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[41] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_97  (.A(
        MAC_MII_COL_net_1), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/COLF_net ), .IPB(), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_246  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[58] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[6] ), .IPC());
    IOINFF_BYPASS \SF2Project_MSS_0/USB_ULPI_DIR_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/USB_ULPI_DIR_PAD_Y ), .Y(
        \SF2Project_MSS_0/USB_ULPI_DIR_PAD/YIN ));
    IOTRI_OB_EB \SF2Project_MSS_0/MDDR_ADDR_11_PAD/U_IOOUT  (.D(VCC), 
        .E(VCC), .DOUT(), .EOUT(
        \SF2Project_MSS_0/MDDR_ADDR_11_PAD/EOUT ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_227  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[11] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[23] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_237  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[35] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[47] ), 
        .IPC());
    sdf_IOPAD_TRI \SF2Project_MSS_0/MDDR_ADDR_11_PAD/U_IOPAD  (.PAD(
        MDDR_ADDR[11]), .D(\SF2Project_MSS_0/DRAM_ADDR_net_0[11] ), .E(
        \SF2Project_MSS_0/MDDR_ADDR_11_PAD/EOUT ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_20  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[25] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_MASTLOCK_net ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_67  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[28] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[1] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_162  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO12A_F2H_GPIN_net ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO15A_F2H_GPIN_net ), .IPC(
        ));
    CFG1 #( .INIT(2'h2) )  BLOCK_INTERFACE_I_MCCC_CLK_BASE (.A(
        MCCC_CLK_BASE), .Y(MCCC_CLK_BASE_net_1));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_7  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[5] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[12] ), .IPC());
    IOBI_IB_OB_EB \SF2Project_MSS_0/MDDR_DQ_11_PAD/U_IOBI  (.D(VCC), 
        .E(VCC), .YIN(\SF2Project_MSS_0/MDDR_DQ_11_PAD/YIN ), .DOUT(), 
        .EOUT(), .Y());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_240  (
        .A(VCC), .B(GND), .C(GND), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[52] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[0] ), .IPC(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WVALID_net ));
    IOINFF_BYPASS \SF2Project_MSS_0/MDDR_DQ_6_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/MDDR_DQ_6_PAD_Y ), .Y(
        \SF2Project_MSS_0/MDDR_DQ_6_PAD/YIN ));
    IOINFF_BYPASS \SF2Project_MSS_0/USB_ULPI_DATA_2_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/USB_ULPI_DATA_2_PAD_Y ), .Y(
        \SF2Project_MSS_0/USB_ULPI_DATA_2_PAD/YIN ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_96  (.A(
        MAC_MII_CRS_net_1), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/CRSF_net ), .IPB(), .IPC());
    sdf_IOPAD_IN \SF2Project_MSS_0/MDDR_DQS_TMATCH_0_IN_PAD/U_IOPAD  (
        .PAD(MDDR_DQS_TMATCH_0_IN), .Y(
        \SF2Project_MSS_0/MDDR_DQS_TMATCH_0_IN_PAD_Y ));
    sdf_IOPAD_TRI \SF2Project_MSS_0/MDDR_ADDR_5_PAD/U_IOPAD  (.PAD(
        MDDR_ADDR[5]), .D(\SF2Project_MSS_0/DRAM_ADDR_net_0[5] ), .E(
        \SF2Project_MSS_0/MDDR_ADDR_5_PAD/EOUT ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_286  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[9] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[13] ), 
        .IPC());
    IO_DIFF \SF2Project_MSS_0/MDDR_DQS_1_PAD/U_ION  (.YIN(GND));
    IOINFF_BYPASS \SF2Project_MSS_0/SPI_1_DI_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/SPI_1_DI_PAD_Y ), .Y(
        \SF2Project_MSS_0/SPI_1_DI_PAD/YIN ));
    IOBI_IB_OB_EB \SF2Project_MSS_0/SPI_1_CLK_PAD/U_IOBI  (.D(VCC), .E(
        VCC), .YIN(\SF2Project_MSS_0/SPI_1_CLK_PAD/YIN ), .DOUT(), 
        .EOUT(), .Y());
    sdf_IOPAD_BI \SF2Project_MSS_0/I2C_1_SCL_PAD/U_IOPAD  (.PAD(
        I2C_1_SCL), .D(
        \SF2Project_MSS_0/MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OUT )
        , .E(
        \SF2Project_MSS_0/MSS_ADLIB_INST_I2C1_SCL_USBA_DATA4_MGPIO1A_OE )
        , .Y(\SF2Project_MSS_0/I2C_1_SCL_PAD_Y ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_208  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[26] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWBURST_HTRANS0_net[0] ), 
        .IPC());
    IOTRI_OB_EB \SF2Project_MSS_0/MDDR_ADDR_6_PAD/U_IOOUT  (.D(VCC), 
        .E(VCC), .DOUT(), .EOUT(
        \SF2Project_MSS_0/MDDR_ADDR_6_PAD/EOUT ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_66  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[27] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[0] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_202  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[6] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[18] )
        , .IPC());
    IOIN_IB \SF2Project_MSS_0/SPI_0_DI_PAD/U_IOIN  (.YIN(
        \SF2Project_MSS_0/SPI_0_DI_PAD/YIN ), .E(GND), .Y());
    IOINFF_BYPASS \SF2Project_MSS_0/USB_ULPI_XCLK_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/USB_ULPI_XCLK_PAD_Y ), .Y(
        \SF2Project_MSS_0/USB_ULPI_XCLK_PAD/YIN ));
    sdf_IOPAD_BI \SF2Project_MSS_0/USB_ULPI_DATA_6_PAD/U_IOPAD  (.PAD(
        USB_ULPI_DATA[6]), .D(
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_TXD3_USBB_DATA6_OUT ), 
        .E(\SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_TXD3_USBB_DATA6_OE ), 
        .Y(\SF2Project_MSS_0/USB_ULPI_DATA_6_PAD_Y ));
    sdf_IOPAD_IN \SF2Project_MSS_0/MMUART_0_RXD_PAD/U_IOPAD  (.PAD(
        MMUART_0_RXD), .Y(\SF2Project_MSS_0/MMUART_0_RXD_PAD_Y ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_225  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[9] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[21] ), 
        .IPC());
    CFG1 #( .INIT(2'h2) )  BLOCK_INTERFACE_I_MAC_MII_TX_CLK (.A(
        MAC_MII_TX_CLK), .Y(MAC_MII_TX_CLK_net_1));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_280  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[3] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[7] ), 
        .IPC());
    sdf_IOPAD_BI \SF2Project_MSS_0/MDDR_DQ_12_PAD/U_IOPAD  (.PAD(
        MDDR_DQ[12]), .D(\SF2Project_MSS_0/DRAM_DQ_OUT_net_0[12] ), .E(
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[12] ), .Y(
        \SF2Project_MSS_0/MDDR_DQ_12_PAD_Y ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_235  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[33] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[45] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_74  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[8] ), 
        .IPB(), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_158  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO10A_F2H_GPIN_net ), .IPB(
        ), .IPC());
    IOINFF_BYPASS \SF2Project_MSS_0/MDDR_DQ_14_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/MDDR_DQ_14_PAD_Y ), .Y(
        \SF2Project_MSS_0/MDDR_DQ_14_PAD/YIN ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_118  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[7] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_141  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2HCALIB_net ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI0_CLK_IN_net ), .IPC());
    IOIN_IB \SF2Project_MSS_0/MDDR_DQS_0_PAD/U_IOP  (.YIN(
        \SF2Project_MSS_0/MDDR_DQS_0_PAD/YIN ), .E(GND), .Y());
    IOIN_IB \SF2Project_MSS_0/USB_ULPI_XCLK_PAD/U_IOIN  (.YIN(
        \SF2Project_MSS_0/USB_ULPI_XCLK_PAD/YIN ), .E(GND), .Y());
    sdf_IOPAD_BI \SF2Project_MSS_0/MDDR_DQ_6_PAD/U_IOPAD  (.PAD(
        MDDR_DQ[6]), .D(\SF2Project_MSS_0/DRAM_DQ_OUT_net_0[6] ), .E(
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[6] ), .Y(
        \SF2Project_MSS_0/MDDR_DQ_6_PAD_Y ));
    IOINFF_BYPASS \SF2Project_MSS_0/MDDR_DQ_4_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/MDDR_DQ_4_PAD_Y ), .Y(
        \SF2Project_MSS_0/MDDR_DQ_4_PAD/YIN ));
    sdf_IOPAD_IN \SF2Project_MSS_0/USB_ULPI_NXT_PAD/U_IOPAD  (.PAD(
        USB_ULPI_NXT), .Y(\SF2Project_MSS_0/USB_ULPI_NXT_PAD_Y ));
    IOINFF_BYPASS \SF2Project_MSS_0/MDDR_DM_RDQS_1_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/MDDR_DM_RDQS_1_PAD_Y ), .Y(
        \SF2Project_MSS_0/MDDR_DM_RDQS_1_PAD/YIN ));
    IOTRI_OB_EB \SF2Project_MSS_0/MDDR_CKE_PAD/U_IOOUT  (.D(VCC), .E(
        VCC), .DOUT(), .EOUT(\SF2Project_MSS_0/MDDR_CKE_PAD/EOUT ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_146  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO0A_F2H_GPIN_net ), .IPB()
        , .IPC());
    sdf_IOPAD_TRI \SF2Project_MSS_0/MDDR_DQS_TMATCH_0_OUT_PAD/U_IOPAD  
        (.PAD(MDDR_DQS_TMATCH_0_OUT), .D(
        \SF2Project_MSS_0/DRAM_FIFO_WE_OUT_net_0[0] ), .E(
        \SF2Project_MSS_0/MDDR_DQS_TMATCH_0_OUT_PAD/EOUT ));
    IOTRI_OB_EB \SF2Project_MSS_0/MDDR_ADDR_15_PAD/U_IOOUT  (.D(VCC), 
        .E(VCC), .DOUT(), .EOUT(
        \SF2Project_MSS_0/MDDR_ADDR_15_PAD/EOUT ));
    sdf_IOPAD_TRI \SF2Project_MSS_0/MDDR_ADDR_13_PAD/U_IOPAD  (.PAD(
        MDDR_ADDR[13]), .D(\SF2Project_MSS_0/DRAM_ADDR_net_0[13] ), .E(
        \SF2Project_MSS_0/MDDR_ADDR_13_PAD/EOUT ));
    sdf_IOPAD_BI \SF2Project_MSS_0/MDDR_DQ_4_PAD/U_IOPAD  (.PAD(
        MDDR_DQ[4]), .D(\SF2Project_MSS_0/DRAM_DQ_OUT_net_0[4] ), .E(
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[4] ), .Y(
        \SF2Project_MSS_0/MDDR_DQ_4_PAD_Y ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_78  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[12] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[19] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_192  (
        .A(GND), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[0] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[8] ), 
        .IPC(\SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[20] )
        );
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_122  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_SESSEND_net ), .IPB(), 
        .IPC());
    sdf_IOPAD_BI \SF2Project_MSS_0/MDDR_DQ_0_PAD/U_IOPAD  (.PAD(
        MDDR_DQ[0]), .D(\SF2Project_MSS_0/DRAM_DQ_OUT_net_0[0] ), .E(
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[0] ), .Y(
        \SF2Project_MSS_0/MDDR_DQ_0_PAD_Y ));
    sdf_IOPAD_TRI \SF2Project_MSS_0/MDDR_BA_1_PAD/U_IOPAD  (.PAD(
        MDDR_BA[1]), .D(\SF2Project_MSS_0/DRAM_BA_net_0[1] ), .E(
        \SF2Project_MSS_0/MDDR_BA_1_PAD/EOUT ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_181  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART0_DCD_F2H_SCP_net ), 
        .IPB(), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_132  (
        .A(GND), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[14] ), .IPB(
        ), .IPC());
    sdf_IOPAD_IN \SF2Project_MSS_0/MMUART_1_RXD_PAD/U_IOPAD  (.PAD(
        MMUART_1_RXD), .Y(\SF2Project_MSS_0/MMUART_1_RXD_PAD_Y ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_45  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[28] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ENABLE_net ), .IPC());
    IOBI_IB_OB_EB \SF2Project_MSS_0/MDDR_DQ_12_PAD/U_IOBI  (.D(VCC), 
        .E(VCC), .YIN(\SF2Project_MSS_0/MDDR_DQ_12_PAD/YIN ), .DOUT(), 
        .EOUT(), .Y());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_99  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/GTX_CLKPF_net ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/RCGF_net[6] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_41  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[24] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[31] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_92  (.A(
        MAC_MII_RX_CLK_net_1), .B(MAC_MII_RX_ER_net_1), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/RX_CLKPF_net ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/RX_ERRF_net ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_2  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[0] ), .IPB(), 
        .IPC());
    IOINFF_BYPASS \SF2Project_MSS_0/I2C_1_SDA_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/I2C_1_SDA_PAD_Y ), .Y(
        \SF2Project_MSS_0/I2C_1_SDA_PAD/YIN ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_93  (.A(
        MAC_MII_RX_DV_net_1), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/RX_DVF_net ), .IPB(), .IPC());
    sdf_IOPAD_TRI \SF2Project_MSS_0/MDDR_ADDR_0_PAD/U_IOPAD  (.PAD(
        MDDR_ADDR[0]), .D(\SF2Project_MSS_0/DRAM_ADDR_net_0[0] ), .E(
        \SF2Project_MSS_0/MDDR_ADDR_0_PAD/EOUT ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_186  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO29B_F2H_GPIN_net ), .IPB(
        ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_178  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART0_DSR_F2H_SCP_net ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_147  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/I2C1_SDA_F2H_SCP_net ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO4A_F2H_GPIN_net ), .IPC()
        );
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_69  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[30] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[3] ), 
        .IPC());
    IOBI_IB_OB_EB \SF2Project_MSS_0/MDDR_DQ_3_PAD/U_IOBI  (.D(VCC), .E(
        VCC), .YIN(\SF2Project_MSS_0/MDDR_DQ_3_PAD/YIN ), .DOUT(), 
        .EOUT(), .Y());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_62  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[23] ), .IPB(), 
        .IPC());
    IOINFF_BYPASS \SF2Project_MSS_0/MDDR_DQS_1_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/MDDR_DQS_1_PAD_Y ), .Y(
        \SF2Project_MSS_0/MDDR_DQS_1_PAD/YIN ));
    sdf_IOPAD_BI \SF2Project_MSS_0/SPI_1_CLK_PAD/U_IOPAD  (.PAD(
        SPI_1_CLK), .D(\SF2Project_MSS_0/MSS_ADLIB_INST_SPI1_SCK_OUT ), 
        .E(\SF2Project_MSS_0/MSS_ADLIB_INST_SPI1_SCK_OE ), .Y(
        \SF2Project_MSS_0/SPI_1_CLK_PAD_Y ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_63  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[24] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[31] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_143  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_M3_RESET_N_net ), .IPC());
    IOBI_IB_OB_EB \SF2Project_MSS_0/I2C_0_SDA_PAD/U_IOBI  (.D(VCC), .E(
        VCC), .YIN(\SF2Project_MSS_0/I2C_0_SDA_PAD/YIN ), .DOUT(), 
        .EOUT(), .Y());
    IOIN_IB \SF2Project_MSS_0/USB_ULPI_NXT_PAD/U_IOIN  (.YIN(
        \SF2Project_MSS_0/USB_ULPI_NXT_PAD/YIN ), .E(GND), .Y());
    IOBI_IB_OB_EB \SF2Project_MSS_0/USB_ULPI_DATA_4_PAD/U_IOBI  (.D(
        VCC), .E(VCC), .YIN(\SF2Project_MSS_0/USB_ULPI_DATA_4_PAD/YIN )
        , .DOUT(), .EOUT(), .Y());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_155  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO8A_F2H_GPIN_net ), .IPC()
        );
    IOTRI_OB_EB \SF2Project_MSS_0/MDDR_ADDR_14_PAD/U_IOOUT  (.D(VCC), 
        .E(VCC), .DOUT(), .EOUT(
        \SF2Project_MSS_0/MDDR_ADDR_14_PAD/EOUT ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_115  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[7] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[4] ), .IPC());
    sdf_IOPAD_TRI \SF2Project_MSS_0/MDDR_ADDR_3_PAD/U_IOPAD  (.PAD(
        MDDR_ADDR[3]), .D(\SF2Project_MSS_0/DRAM_ADDR_net_0[3] ), .E(
        \SF2Project_MSS_0/MDDR_ADDR_3_PAD/EOUT ));
    IOTRI_OB_EB \SF2Project_MSS_0/MDDR_ADDR_12_PAD/U_IOOUT  (.D(VCC), 
        .E(VCC), .DOUT(), .EOUT(
        \SF2Project_MSS_0/MDDR_ADDR_12_PAD/EOUT ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_168  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART1_CTS_F2H_SCP_net ), 
        .IPB(), .IPC());
    sdf_IOPAD_BI \SF2Project_MSS_0/MDDR_DQ_1_PAD/U_IOPAD  (.PAD(
        MDDR_DQ[1]), .D(\SF2Project_MSS_0/DRAM_DQ_OUT_net_0[1] ), .E(
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[1] ), .Y(
        \SF2Project_MSS_0/MDDR_DQ_1_PAD_Y ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_187  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART0_SCK_F2H_SCP_net ), 
        .IPB(), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_24  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[0] ), .IPB(), 
        .IPC());
    IOBI_IB_OB_EB \SF2Project_MSS_0/MDDR_DQ_9_PAD/U_IOBI  (.D(VCC), .E(
        VCC), .YIN(\SF2Project_MSS_0/MDDR_DQ_9_PAD/YIN ), .DOUT(), 
        .EOUT(), .Y());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_47  (.A(
        VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[1] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_183  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART0_TXD_F2H_SCP_net ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/MMUART0_RI_F2H_SCP_net ), 
        .IPC());
    IOTRI_OB_EB \SF2Project_MSS_0/MDDR_ADDR_1_PAD/U_IOOUT  (.D(VCC), 
        .E(VCC), .DOUT(), .EOUT(
        \SF2Project_MSS_0/MDDR_ADDR_1_PAD/EOUT ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_209  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[27] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWBURST_HTRANS0_net[1] ), 
        .IPC());
    CFG1 #( .INIT(2'h2) )  \BLOCK_INTERFACE_I_MAC_MII_RXD[0]  (.A(
        MAC_MII_RXD[0]), .Y(\MAC_MII_RXD[0] ));
    IOINFF_BYPASS \SF2Project_MSS_0/MDDR_DQ_5_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/MDDR_DQ_5_PAD_Y ), .Y(
        \SF2Project_MSS_0/MDDR_DQ_5_PAD/YIN ));
    IOINFF_BYPASS \SF2Project_MSS_0/I2C_0_SDA_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/I2C_0_SDA_PAD_Y ), .Y(
        \SF2Project_MSS_0/I2C_0_SDA_PAD/YIN ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_10  (.A(
        VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[15] ), .IPC());
    IOIN_IB \SF2Project_MSS_0/MMUART_0_RXD_PAD/U_IOIN  (.YIN(
        \SF2Project_MSS_0/MMUART_0_RXD_PAD/YIN ), .E(GND), .Y());
    IOBI_IB_OB_EB \SF2Project_MSS_0/USB_ULPI_DATA_0_PAD/U_IOBI  (.D(
        VCC), .E(VCC), .YIN(\SF2Project_MSS_0/USB_ULPI_DATA_0_PAD/YIN )
        , .DOUT(), .EOUT(), .Y());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_248  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[60] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[0] ), 
        .IPC());
    IOTRI_OB_EB \SF2Project_MSS_0/MDDR_ADDR_2_PAD/U_IOOUT  (.D(VCC), 
        .E(VCC), .DOUT(), .EOUT(
        \SF2Project_MSS_0/MDDR_ADDR_2_PAD/EOUT ));
    CFG1 #( .INIT(2'h2) )  BLOCK_INTERFACE_I_MAC_MII_COL (.A(
        MAC_MII_COL), .Y(MAC_MII_COL_net_1));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_28  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[4] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[11] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_242  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[54] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[2] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_46  (.A(
        VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[0] ), .IPC());
    IOTRI_OB_EB \SF2Project_MSS_0/MMUART_0_TXD_PAD/U_IOOUT  (.D(VCC), 
        .E(VCC), .DOUT(), .EOUT());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_175  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART1_SCK_F2H_SCP_net ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO19B_F2H_GPIN_net ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_204  (
        .A(VCC), .B(GND), .C(GND), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[22] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[0] ), 
        .IPC(\SF2Project_MSS_0/MSS_ADLIB_INST/F_AWVALID_HWRITE0_net ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_104  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/RCGF_net[4] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_LINESTATE_net[0] ), .IPC()
        );
    IOBI_IB_OB_EB \SF2Project_MSS_0/MDDR_DQ_1_PAD/U_IOBI  (.D(VCC), .E(
        VCC), .YIN(\SF2Project_MSS_0/MDDR_DQ_1_PAD/YIN ), .DOUT(), 
        .EOUT(), .Y());
    IO_DIFF \SF2Project_MSS_0/MDDR_CLK_PAD/U_IOP  (.YIN(GND));
    sdf_IOPAD_TRI \SF2Project_MSS_0/MDDR_ADDR_14_PAD/U_IOPAD  (.PAD(
        MDDR_ADDR[14]), .D(\SF2Project_MSS_0/DRAM_ADDR_net_0[14] ), .E(
        \SF2Project_MSS_0/MDDR_ADDR_14_PAD/EOUT ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_50  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[4] ), .IPB(), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_256  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[4] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[16] )
        , .IPC());
    CFG1 #( .INIT(2'h2) )  \BLOCK_INTERFACE_I_MAC_MII_RXD[1]  (.A(
        MAC_MII_RXD[1]), .Y(\MAC_MII_RXD[1] ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_216  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[0] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[12] ), 
        .IPC(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[24] ));
    sdf_IOPAD_BI \SF2Project_MSS_0/MDDR_DM_RDQS_0_PAD/U_IOPAD  (.PAD(
        MDDR_DM_RDQS[0]), .D(
        \SF2Project_MSS_0/DRAM_DM_RDQS_OUT_net_0[0] ), .E(
        \SF2Project_MSS_0/DM_OE_net_0[0] ), .Y(
        \SF2Project_MSS_0/MDDR_DM_RDQS_0_PAD_Y ));
    sdf_IOPAD_BI \SF2Project_MSS_0/USB_ULPI_DATA_1_PAD/U_IOPAD  (.PAD(
        USB_ULPI_DATA[1]), .D(
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT )
        , .E(
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE )
        , .Y(\SF2Project_MSS_0/USB_ULPI_DATA_1_PAD_Y ));
    IOBI_IB_OB_EB \SF2Project_MSS_0/SPI_0_SS0_PAD/U_IOBI  (.D(VCC), .E(
        VCC), .YIN(\SF2Project_MSS_0/SPI_0_SS0_PAD/YIN ), .DOUT(), 
        .EOUT(), .Y());
    IOTRI_OB_EB \SF2Project_MSS_0/MDDR_ADDR_0_PAD/U_IOOUT  (.D(VCC), 
        .E(VCC), .DOUT(), .EOUT(
        \SF2Project_MSS_0/MDDR_ADDR_0_PAD/EOUT ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_109  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[1] ), .IPB(), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_30  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[6] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[13] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_282  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[5] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[9] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_165  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI1_SS0_F2H_SCP_net ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI1_SS3_F2H_SCP_net ), .IPC()
        );
    IOINFF_BYPASS \SF2Project_MSS_0/MDDR_DQ_3_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/MDDR_DQ_3_PAD_Y ), .Y(
        \SF2Project_MSS_0/MDDR_DQ_3_PAD/YIN ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_100  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/RCGF_net[0] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/RCGF_net[7] ), .IPC());
    sdf_IOPAD_BI \SF2Project_MSS_0/USB_ULPI_DATA_5_PAD/U_IOPAD  (.PAD(
        USB_ULPI_DATA[5]), .D(
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_TXD2_USBB_DATA5_OUT ), 
        .E(\SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_TXD2_USBB_DATA5_OE ), 
        .Y(\SF2Project_MSS_0/USB_ULPI_DATA_5_PAD_Y ));
    IOBI_IB_OB_EB \SF2Project_MSS_0/MDDR_DQ_4_PAD/U_IOBI  (.D(VCC), .E(
        VCC), .YIN(\SF2Project_MSS_0/MDDR_DQ_4_PAD/YIN ), .DOUT(), 
        .EOUT(), .Y());
    sdf_IOPAD_TRI \SF2Project_MSS_0/SPI_0_DO_PAD/U_IOPAD  (.PAD(
        SPI_0_DO), .D(
        \SF2Project_MSS_0/MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OUT )
        , .E(
        \SF2Project_MSS_0/MSS_ADLIB_INST_SPI0_SDO_USBA_STP_MGPIO6A_OE )
        );
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_250  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[62] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[2] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_210  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[28] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWLOCK_HMASTLOCK0_net[0] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_198  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[2] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[14] )
        , .IPC());
    IOINFF_BYPASS \SF2Project_MSS_0/SPI_0_DI_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/SPI_0_DI_PAD_Y ), .Y(
        \SF2Project_MSS_0/SPI_0_DI_PAD/YIN ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_128  (
        .A(GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[3] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[10] ), .IPC(
        ));
    sdf_IOPAD_BI \SF2Project_MSS_0/MDDR_DQ_8_PAD/U_IOPAD  (.PAD(
        MDDR_DQ[8]), .D(\SF2Project_MSS_0/DRAM_DQ_OUT_net_0[8] ), .E(
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[8] ), .Y(
        \SF2Project_MSS_0/MDDR_DQ_8_PAD_Y ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_138  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/SMBALERT_NI1_net ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2_DMAREADY_net[0] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_80  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[14] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[21] ), 
        .IPC());
    IOTRI_OB_EB \SF2Project_MSS_0/MDDR_ADDR_5_PAD/U_IOOUT  (.D(VCC), 
        .E(VCC), .DOUT(), .EOUT(
        \SF2Project_MSS_0/MDDR_ADDR_5_PAD/EOUT ));
    CFG1 #( .INIT(2'h2) )  BLOCK_INTERFACE_I_MAC_MII_TX_EN (.A(
        MAC_MII_TX_EN_net_1), .Y(MAC_MII_TX_EN));
    IOTRI_OB_EB \SF2Project_MSS_0/SPI_1_DO_PAD/U_IOOUT  (.D(VCC), .E(
        VCC), .DOUT(), .EOUT());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_276  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[0] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[3] ), 
        .IPC(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[15] ));
    IOBI_IB_OB_EB \SF2Project_MSS_0/MDDR_DQ_10_PAD/U_IOBI  (.D(VCC), 
        .E(VCC), .YIN(\SF2Project_MSS_0/MDDR_DQ_10_PAD/YIN ), .DOUT(), 
        .EOUT(), .Y());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_75  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[9] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[16] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_49  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[3] ), .IPB(), 
        .IPC());
    IOINFF_BYPASS \SF2Project_MSS_0/SPI_1_SS0_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/SPI_1_SS0_PAD_Y ), .Y(
        \SF2Project_MSS_0/SPI_1_SS0_PAD/YIN ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_71  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[5] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_42  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[25] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WRITE_net ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_1  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RESP_net ), .IPB(), 
        .IPC());
    sdf_IOPAD_BI \SF2Project_MSS_0/MDDR_DQ_14_PAD/U_IOPAD  (.PAD(
        MDDR_DQ[14]), .D(\SF2Project_MSS_0/DRAM_DQ_OUT_net_0[14] ), .E(
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[14] ), .Y(
        \SF2Project_MSS_0/MDDR_DQ_14_PAD_Y ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_43  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[26] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_SEL_net ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_151  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/CAN_TXBUS_F2H_SCP_net ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO6A_F2H_GPIN_net ), .IPC()
        );
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_111  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[3] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[0] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_270  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[30] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_RREADY_net ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_266  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[26] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARLOCK_HMASTLOCK1_net[0] ), 
        .IPC());
    IOTRI_OB_EB \SF2Project_MSS_0/MDDR_ADDR_10_PAD/U_IOOUT  (.D(VCC), 
        .E(VCC), .DOUT(), .EOUT(
        \SF2Project_MSS_0/MDDR_ADDR_10_PAD/EOUT ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_156  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO9A_F2H_GPIN_net ), .IPB()
        , .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_116  (
        .A(GND), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_RXVALIDH_net ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[5] ), .IPC());
    IOINFF_BYPASS \SF2Project_MSS_0/MDDR_DQ_2_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/MDDR_DQ_2_PAD_Y ), .Y(
        \SF2Project_MSS_0/MDDR_DQ_2_PAD/YIN ));
    IOINFF_BYPASS \SF2Project_MSS_0/SPI_0_CLK_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/SPI_0_CLK_PAD_Y ), .Y(
        \SF2Project_MSS_0/SPI_0_CLK_PAD/YIN ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_5  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[3] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[10] ), .IPC());
    sdf_IOPAD_TRI \SF2Project_MSS_0/MMUART_1_TXD_PAD/U_IOPAD  (.PAD(
        MMUART_1_TXD), .D(
        \SF2Project_MSS_0/MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT )
        , .E(
        \SF2Project_MSS_0/MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OE )
        );
    IO_DIFF \SF2Project_MSS_0/MDDR_DQS_0_PAD/U_ION  (.YIN(GND));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_195  (
        .A(GND), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[3] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[11] ), 
        .IPC());
    IOBI_IB_OB_EB \SF2Project_MSS_0/MDDR_DM_RDQS_0_PAD/U_IOBI  (.D(VCC)
        , .E(VCC), .YIN(\SF2Project_MSS_0/MDDR_DM_RDQS_0_PAD/YIN ), 
        .DOUT(), .EOUT(), .Y());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_203  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[7] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[19] )
        , .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_125  (
        .A(GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[0] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[7] ), .IPC()
        );
    sdf_IOPAD_BI \SF2Project_MSS_0/I2C_1_SDA_PAD/U_IOPAD  (.PAD(
        I2C_1_SDA), .D(
        \SF2Project_MSS_0/MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OUT )
        , .E(
        \SF2Project_MSS_0/MSS_ADLIB_INST_I2C1_SDA_USBA_DATA3_MGPIO0A_OE )
        , .Y(\SF2Project_MSS_0/I2C_1_SDA_PAD_Y ));
    CFG1 #( .INIT(2'h2) )  BLOCK_INTERFACE_I_MAC_MII_RX_ER (.A(
        MAC_MII_RX_ER), .Y(MAC_MII_RX_ER_net_1));
    IOINFF_BYPASS \SF2Project_MSS_0/USB_ULPI_DATA_0_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/USB_ULPI_DATA_0_PAD_Y ), .Y(
        \SF2Project_MSS_0/USB_ULPI_DATA_0_PAD/YIN ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_260  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[8] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[20] )
        , .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_249  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[61] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[1] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_201  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[5] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[17] )
        , .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_135  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/SMBALERT_NI0_net ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/USER_MSS_RESET_N_net ), .IPC()
        );
    sdf_IOPAD_TRI \SF2Project_MSS_0/MDDR_RESET_N_PAD/U_IOPAD  (.PAD(
        MDDR_RESET_N), .D(\SF2Project_MSS_0/MSS_ADLIB_INST_DRAM_RSTN ), 
        .E(\SF2Project_MSS_0/MDDR_RESET_N_PAD/EOUT ));
    IOTRI_OB_EB \SF2Project_MSS_0/MDDR_ADDR_7_PAD/U_IOOUT  (.D(VCC), 
        .E(VCC), .DOUT(), .EOUT(
        \SF2Project_MSS_0/MDDR_ADDR_7_PAD/EOUT ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_3  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[1] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[8] ), .IPC());
    sdf_IOPAD_TRI \SF2Project_MSS_0/MDDR_ADDR_15_PAD/U_IOPAD  (.PAD(
        MDDR_ADDR[15]), .D(\SF2Project_MSS_0/DRAM_ADDR_net_0[15] ), .E(
        \SF2Project_MSS_0/MDDR_ADDR_15_PAD/EOUT ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_14  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[19] ), .IPB(), 
        .IPC());
    IOBI_IB_OB_EB \SF2Project_MSS_0/MDDR_DQ_2_PAD/U_IOBI  (.D(VCC), .E(
        VCC), .YIN(\SF2Project_MSS_0/MDDR_DQ_2_PAD/YIN ), .DOUT(), 
        .EOUT(), .Y());
    sdf_IOPAD_IN \SF2Project_MSS_0/USB_ULPI_DIR_PAD/U_IOPAD  (.PAD(
        USB_ULPI_DIR), .Y(\SF2Project_MSS_0/USB_ULPI_DIR_PAD_Y ));
    sdf_IOPAD_IN \SF2Project_MSS_0/SPI_1_DI_PAD/U_IOPAD  (.PAD(
        SPI_1_DI), .Y(\SF2Project_MSS_0/SPI_1_DI_PAD_Y ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_77  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[11] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[18] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_207  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[25] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[3] ), 
        .IPC());
    IOBI_IB_OB_EB \SF2Project_MSS_0/MDDR_DM_RDQS_1_PAD/U_IOBI  (.D(VCC)
        , .E(VCC), .YIN(\SF2Project_MSS_0/MDDR_DM_RDQS_1_PAD/YIN ), 
        .DOUT(), .EOUT(), .Y());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_157  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI0_SS2_F2H_SCP_net ), .IPB()
        , .IPC());
    sdf_IOPAD_TRI \SF2Project_MSS_0/MDDR_ADDR_4_PAD/U_IOPAD  (.PAD(
        MDDR_ADDR[4]), .D(\SF2Project_MSS_0/DRAM_ADDR_net_0[4] ), .E(
        \SF2Project_MSS_0/MDDR_ADDR_4_PAD/EOUT ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_117  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_RXACTIVE_net ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[6] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_171  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART1_DCD_F2H_SCP_net ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO17B_F2H_GPIN_net ), 
        .IPC());
    sdf_IOPAD_TRI \SF2Project_MSS_0/MDDR_WE_N_PAD/U_IOPAD  (.PAD(
        MDDR_WE_N), .D(\SF2Project_MSS_0/MSS_ADLIB_INST_DRAM_WEN ), .E(
        \SF2Project_MSS_0/MDDR_WE_N_PAD/EOUT ));
    sdf_IOPAD_BI \SF2Project_MSS_0/MDDR_DM_RDQS_1_PAD/U_IOPAD  (.PAD(
        MDDR_DM_RDQS[1]), .D(
        \SF2Project_MSS_0/DRAM_DM_RDQS_OUT_net_0[1] ), .E(
        \SF2Project_MSS_0/DM_OE_net_0[1] ), .Y(
        \SF2Project_MSS_0/MDDR_DM_RDQS_1_PAD_Y ));
    sdf_IOPAD_TRI \SF2Project_MSS_0/MDDR_ADDR_7_PAD/U_IOPAD  (.PAD(
        MDDR_ADDR[7]), .D(\SF2Project_MSS_0/DRAM_ADDR_net_0[7] ), .E(
        \SF2Project_MSS_0/MDDR_ADDR_7_PAD/EOUT ));
    IOINFF_BYPASS \SF2Project_MSS_0/MDDR_DQ_10_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/MDDR_DQ_10_PAD_Y ), .Y(
        \SF2Project_MSS_0/MDDR_DQ_10_PAD/YIN ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_153  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/CAN_RXBUS_F2H_SCP_net ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO7A_F2H_GPIN_net ), .IPC()
        );
    sdf_IOPAD_TRI \SF2Project_MSS_0/MMUART_0_TXD_PAD/U_IOPAD  (.PAD(
        MMUART_0_TXD), .D(
        \SF2Project_MSS_0/MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OUT )
        , .E(
        \SF2Project_MSS_0/MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OE )
        );
    IOINFF_BYPASS \SF2Project_MSS_0/USB_ULPI_DATA_6_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/USB_ULPI_DATA_6_PAD_Y ), .Y(
        \SF2Project_MSS_0/USB_ULPI_DATA_6_PAD/YIN ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_8  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[6] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[13] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_113  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[5] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[2] ), .IPC());
    CFG1 #( .INIT(2'h2) )  \BLOCK_INTERFACE_I_MAC_MII_RXD[2]  (.A(
        MAC_MII_RXD[2]), .Y(\MAC_MII_RXD[2] ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_244  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[56] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[4] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_144  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_PLL_LOCK_net ), .IPB(), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_54  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[8] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[15] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_18  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[23] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[30] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_176  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO26B_F2H_GPIN_net ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART0_CTS_F2H_SCP_net ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_76  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[10] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[17] ), 
        .IPC());
    sdf_IOPAD_BI \SF2Project_MSS_0/MDDR_DQ_10_PAD/U_IOPAD  (.PAD(
        MDDR_DQ[10]), .D(\SF2Project_MSS_0/DRAM_DQ_OUT_net_0[10] ), .E(
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[10] ), .Y(
        \SF2Project_MSS_0/MDDR_DQ_10_PAD_Y ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_149  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/I2C1_SCL_F2H_SCP_net ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO5A_F2H_GPIN_net ), .IPC()
        );
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_34  (.A(
        VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[17] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_161  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI1_SDI_F2H_SCP_net ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI1_SS1_F2H_SCP_net ), .IPC()
        );
    IOINFF_BYPASS \SF2Project_MSS_0/MDDR_DQ_7_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/MDDR_DQ_7_PAD_Y ), .Y(
        \SF2Project_MSS_0/MDDR_DQ_7_PAD/YIN ));
    sdf_IOPAD_TRI \SF2Project_MSS_0/MDDR_CKE_PAD/U_IOPAD  (.PAD(
        MDDR_CKE), .D(\SF2Project_MSS_0/MSS_ADLIB_INST_DRAM_CKE ), .E(
        \SF2Project_MSS_0/MDDR_CKE_PAD/EOUT ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_25  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[1] ), .IPB(), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_21  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[26] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_SIZE_net[0] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_140  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/RX_EV_net ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/USER_MSS_GPIO_RESET_N_net ), 
        .IPC());
    IOBI_IB_OB_EB \SF2Project_MSS_0/MDDR_DQ_15_PAD/U_IOBI  (.D(VCC), 
        .E(VCC), .YIN(\SF2Project_MSS_0/MDDR_DQ_15_PAD/YIN ), .DOUT(), 
        .EOUT(), .Y());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_226  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[10] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[22] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_205  (
        .A(VCC), .B(GND), .C(GND), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[23] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[1] ), 
        .IPC(\SF2Project_MSS_0/MSS_ADLIB_INST/F_WLAST_net ));
    CFG1 #( .INIT(2'h2) )  BLOCK_INTERFACE_I_MAC_MII_TX_ER (.A(
        MAC_MII_TX_ER_net_1), .Y(MAC_MII_TX_ER));
    CFG1 #( .INIT(2'h2) )  \BLOCK_INTERFACE_I_MAC_MII_RXD[3]  (.A(
        MAC_MII_RXD[3]), .Y(\MAC_MII_RXD[3] ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_284  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[7] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[11] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_236  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[34] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[46] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_184  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO28B_F2H_GPIN_net ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO31B_F2H_GPIN_net ), .IPC(
        ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_58  (.A(
        VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[19] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_166  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO11B_F2H_GPIN_net ), .IPC(
        ));
    sdf_IOPAD_TRI \SF2Project_MSS_0/MDDR_CS_N_PAD/U_IOPAD  (.PAD(
        MDDR_CS_N), .D(\SF2Project_MSS_0/MSS_ADLIB_INST_DRAM_CSN ), .E(
        \SF2Project_MSS_0/MDDR_CS_N_PAD/EOUT ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_177  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART1_RXD_F2H_SCP_net ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO20B_F2H_GPIN_net ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_84  (.A(
        VCC), .B(\MAC_MII_RXD[0] ), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[25] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/RXDF_net[0] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_258  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[6] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[18] )
        , .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_189  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/I2C0_SDA_F2H_SCP_net ), .IPB()
        , .IPC());
    IOINFF_BYPASS \SF2Project_MSS_0/I2C_0_SCL_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/I2C_0_SCL_PAD_Y ), .Y(
        \SF2Project_MSS_0/I2C_0_SCL_PAD/YIN ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_38  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[21] ), .IPB(), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_218  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[2] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[14] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_173  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART1_TXD_F2H_SCP_net ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO18B_F2H_GPIN_net ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_252  (
        .A(VCC), .B(VCC), .C(GND), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[0] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[12] )
        , .IPC(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARSIZE_HSIZE1_net[0] ));
    sdf_IOPAD_BI \SF2Project_MSS_0/USB_ULPI_DATA_4_PAD/U_IOPAD  (.PAD(
        USB_ULPI_DATA[4]), .D(
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_RXD3_USBB_DATA4_OUT ), 
        .E(\SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_RXD3_USBB_DATA4_OE ), 
        .Y(\SF2Project_MSS_0/USB_ULPI_DATA_4_PAD_Y ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_220  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[4] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[16] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_212  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[30] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[0] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_230  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[28] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[40] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_180  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO22B_F2H_GPIN_net ), .IPB(
        ), .IPC());
    IOIN_IB \SF2Project_MSS_0/MMUART_1_RXD_PAD/U_IOIN  (.YIN(
        \SF2Project_MSS_0/MMUART_1_RXD_PAD/YIN ), .E(GND), .Y());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_167  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MMUART1_RTS_F2H_SCP_net ), 
        .IPC());
    IOINFF_BYPASS \SF2Project_MSS_0/MDDR_DQ_1_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/MDDR_DQ_1_PAD_Y ), .Y(
        \SF2Project_MSS_0/MDDR_DQ_1_PAD/YIN ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_88  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[29] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/RXDF_net[4] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_27  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[3] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[10] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_163  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI1_SDO_F2H_SCP_net ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI1_SS2_F2H_SCP_net ), .IPC()
        );
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_102  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/RCGF_net[2] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/RCGF_net[9] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_90  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[31] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/RXDF_net[6] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_79  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[13] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[20] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_72  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[6] ), 
        .IPB(), .IPC());
    sdf_IOPAD_BI \SF2Project_MSS_0/USB_ULPI_DATA_3_PAD/U_IOPAD  (.PAD(
        USB_ULPI_DATA[3]), .D(
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT )
        , .E(
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE )
        , .Y(\SF2Project_MSS_0/USB_ULPI_DATA_3_PAD_Y ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_73  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[7] ), 
        .IPB(), .IPC());
    IOINFF_BYPASS \SF2Project_MSS_0/MMUART_0_RXD_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/MMUART_0_RXD_PAD_Y ), .Y(
        \SF2Project_MSS_0/MMUART_0_RXD_PAD/YIN ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_278  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[2] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[5] ), 
        .IPC());
    IOTRI_OB_EB \SF2Project_MSS_0/MMUART_1_TXD_PAD/U_IOOUT  (.D(VCC), 
        .E(VCC), .DOUT(), .EOUT());
    IOTRI_OB_EB \SF2Project_MSS_0/MDDR_WE_N_PAD/U_IOOUT  (.D(VCC), .E(
        VCC), .DOUT(), .EOUT(\SF2Project_MSS_0/MDDR_WE_N_PAD/EOUT ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_26  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[2] ), .IPB(), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_121  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_AVALID_net ), .IPB(), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_60  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[21] ), .IPB(), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_272  (
        .A(GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[0] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_RMW_AXI_net ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_131  (
        .A(VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[13] ), .IPC(
        ));
    IOTRI_OB_EB \SF2Project_MSS_0/MDDR_ODT_PAD/U_IOOUT  (.D(VCC), .E(
        VCC), .DOUT(), .EOUT(\SF2Project_MSS_0/MDDR_ODT_PAD/EOUT ));
    sdf_IOPAD_TRI \SF2Project_MSS_0/MDDR_ADDR_6_PAD/U_IOPAD  (.PAD(
        MDDR_ADDR[6]), .D(\SF2Project_MSS_0/DRAM_ADDR_net_0[6] ), .E(
        \SF2Project_MSS_0/MDDR_ADDR_6_PAD/EOUT ));
    IOBI_IB_OB_EB \SF2Project_MSS_0/USB_ULPI_DATA_7_PAD/U_IOBI  (.D(
        VCC), .E(VCC), .YIN(\SF2Project_MSS_0/USB_ULPI_DATA_7_PAD/YIN )
        , .DOUT(), .EOUT(), .Y());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_243  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[55] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[3] ), .IPC());
    IOBI_IB_OB_EB \SF2Project_MSS_0/SPI_0_CLK_PAD/U_IOBI  (.D(VCC), .E(
        VCC), .YIN(\SF2Project_MSS_0/SPI_0_CLK_PAD/YIN ), .DOUT(), 
        .EOUT(), .Y());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_241  (
        .A(VCC), .B(GND), .C(GND), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[53] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[1] ), .IPC(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_BREADY_net ));
    IOBI_IB_OB_EB \SF2Project_MSS_0/MDDR_DQ_0_PAD/U_IOBI  (.D(VCC), .E(
        VCC), .YIN(\SF2Project_MSS_0/MDDR_DQ_0_PAD/YIN ), .DOUT(), 
        .EOUT(), .Y());
    IOINFF_BYPASS \SF2Project_MSS_0/SPI_1_CLK_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/SPI_1_CLK_PAD_Y ), .Y(
        \SF2Project_MSS_0/SPI_1_CLK_PAD/YIN ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_196  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[0] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[12] )
        , .IPC());
    sdf_IOPAD_TRI \SF2Project_MSS_0/MDDR_BA_2_PAD/U_IOPAD  (.PAD(
        MDDR_BA[2]), .D(\SF2Project_MSS_0/DRAM_BA_net_0[2] ), .E(
        \SF2Project_MSS_0/MDDR_BA_2_PAD/EOUT ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_126  (
        .A(GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[1] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[8] ), .IPC()
        );
    IOTRI_OB_EB \SF2Project_MSS_0/MDDR_CAS_N_PAD/U_IOOUT  (.D(VCC), .E(
        VCC), .DOUT(), .EOUT(\SF2Project_MSS_0/MDDR_CAS_N_PAD/EOUT ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_136  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/SMBSUS_NI0_net ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_DMAREADY_net[0] ), .IPC());
    IOIN_IB \SF2Project_MSS_0/MDDR_DQS_TMATCH_0_IN_PAD/U_IOIN  (.YIN(
        \SF2Project_MSS_0/MDDR_DQS_TMATCH_0_IN_PAD/YIN ), .E(GND), .Y()
        );
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_247  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[59] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[7] ), .IPC());
    IOIN_IB \SF2Project_MSS_0/SPI_1_DI_PAD/U_IOIN  (.YIN(
        \SF2Project_MSS_0/SPI_1_DI_PAD/YIN ), .E(GND), .Y());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_268  (
        .A(VCC), .B(MCCC_CLK_BASE_net_1), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[28] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/CLK_BASE_net ), .IPC());
    IOBI_IB_OB_EB \SF2Project_MSS_0/I2C_1_SCL_PAD/U_IOBI  (.D(VCC), .E(
        VCC), .YIN(\SF2Project_MSS_0/I2C_1_SCL_PAD/YIN ), .DOUT(), 
        .EOUT(), .Y());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_262  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[10] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[22] )
        , .IPC());
    IOBI_IB_OB_EB \SF2Project_MSS_0/MDDR_DQ_7_PAD/U_IOBI  (.D(VCC), .E(
        VCC), .YIN(\SF2Project_MSS_0/MDDR_DQ_7_PAD/YIN ), .DOUT(), 
        .EOUT(), .Y());
    IOTRI_OB_EB \SF2Project_MSS_0/MDDR_ADDR_4_PAD/U_IOOUT  (.D(VCC), 
        .E(VCC), .DOUT(), .EOUT(
        \SF2Project_MSS_0/MDDR_ADDR_4_PAD/EOUT ));
    IOINFF_BYPASS \SF2Project_MSS_0/MDDR_DQ_8_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/MDDR_DQ_8_PAD_Y ), .Y(
        \SF2Project_MSS_0/MDDR_DQ_8_PAD/YIN ));
    IOINFF_BYPASS \SF2Project_MSS_0/MDDR_DQ_15_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/MDDR_DQ_15_PAD_Y ), .Y(
        \SF2Project_MSS_0/MDDR_DQ_15_PAD/YIN ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_283  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[6] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[10] ), 
        .IPC());
    IOINFF_BYPASS \SF2Project_MSS_0/USB_ULPI_NXT_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/USB_ULPI_NXT_PAD_Y ), .Y(
        \SF2Project_MSS_0/USB_ULPI_NXT_PAD/YIN ));
    sdf_IOPAD_BI \SF2Project_MSS_0/USB_ULPI_DATA_7_PAD/U_IOPAD  (.PAD(
        USB_ULPI_DATA[7]), .D(
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT )
        , .E(
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE )
        , .Y(\SF2Project_MSS_0/USB_ULPI_DATA_7_PAD_Y ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_281  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[4] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[8] ), 
        .IPC());
    sdf_IOPAD_BI \SF2Project_MSS_0/MDDR_DQ_15_PAD/U_IOPAD  (.PAD(
        MDDR_DQ[15]), .D(\SF2Project_MSS_0/DRAM_DQ_OUT_net_0[15] ), .E(
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[15] ), .Y(
        \SF2Project_MSS_0/MDDR_DQ_15_PAD_Y ));
    IOTRI_OB_EB \SF2Project_MSS_0/MDDR_RAS_N_PAD/U_IOOUT  (.D(VCC), .E(
        VCC), .DOUT(), .EOUT(\SF2Project_MSS_0/MDDR_RAS_N_PAD/EOUT ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_197  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[1] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[13] )
        , .IPC());
    sdf_IOPAD_TRI \SF2Project_MSS_0/MDDR_ODT_PAD/U_IOPAD  (.PAD(
        MDDR_ODT), .D(\SF2Project_MSS_0/MSS_ADLIB_INST_DRAM_ODT ), .E(
        \SF2Project_MSS_0/MDDR_ODT_PAD/EOUT ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_127  (
        .A(GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[2] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[9] ), .IPC()
        );
    sdf_IOPADP_BI \SF2Project_MSS_0/MDDR_DQS_1_PAD/U_IOPADP  (.PAD_P(
        MDDR_DQS[1]), .N2PIN_P(
        \SF2Project_MSS_0/MDDR_DQS_1_PAD/U2_N2P ), .OIN_P(
        \SF2Project_MSS_0/DRAM_DQS_OUT_net_0[1] ), .EIN_P(
        \SF2Project_MSS_0/DRAM_DQS_OE_net_0[1] ), .IOUT_P(
        \SF2Project_MSS_0/MDDR_DQS_1_PAD_Y ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_287  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[10] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[14] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_137  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/I2C1_BCLK_net ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_DMAREADY_net[1] ), .IPC());
    sdf_IOPAD_TRI \SF2Project_MSS_0/USB_ULPI_STP_PAD/U_IOPAD  (.PAD(
        USB_ULPI_STP), .D(
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_TXD1_RMII_TXD1_USBB_STP_OUT )
        , .E(
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_TXD1_RMII_TXD1_USBB_STP_OE )
        );
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_193  (
        .A(GND), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[1] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[9] ), 
        .IPC(\SF2Project_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[21] )
        );
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_123  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_HOSTDISCON_net ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[5] ), .IPC()
        );
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_133  (
        .A(GND), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[15] ), .IPB(
        ), .IPC());
    sdf_IOPAD_BI \SF2Project_MSS_0/SPI_1_SS0_PAD/U_IOPAD  (.PAD(
        SPI_1_SS0), .D(
        \SF2Project_MSS_0/MSS_ADLIB_INST_SPI1_SS0_MGPIO13A_OUT ), .E(
        \SF2Project_MSS_0/MSS_ADLIB_INST_SPI1_SS0_MGPIO13A_OE ), .Y(
        \SF2Project_MSS_0/SPI_1_SS0_PAD_Y ));
    sdf_IOPAD_BI \SF2Project_MSS_0/MDDR_DQ_7_PAD/U_IOPAD  (.PAD(
        MDDR_DQ[7]), .D(\SF2Project_MSS_0/DRAM_DQ_OUT_net_0[7] ), .E(
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[7] ), .Y(
        \SF2Project_MSS_0/MDDR_DQ_7_PAD_Y ));
    IOINFF_BYPASS \SF2Project_MSS_0/MDDR_DQS_0_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/MDDR_DQS_0_PAD_Y ), .Y(
        \SF2Project_MSS_0/MDDR_DQS_0_PAD/YIN ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_245  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[57] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[5] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_259  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[7] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[19] )
        , .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_219  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[3] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[15] ), 
        .IPC());
    sdf_IOPAD_BI \SF2Project_MSS_0/MDDR_DQ_9_PAD/U_IOPAD  (.PAD(
        MDDR_DQ[9]), .D(\SF2Project_MSS_0/DRAM_DQ_OUT_net_0[9] ), .E(
        \SF2Project_MSS_0/DRAM_DQ_OE_net_0[9] ), .Y(
        \SF2Project_MSS_0/MDDR_DQ_9_PAD_Y ));
    IOINFF_BYPASS \SF2Project_MSS_0/MDDR_DQS_TMATCH_0_IN_PAD/U_IOINFF  
        (.A(\SF2Project_MSS_0/MDDR_DQS_TMATCH_0_IN_PAD_Y ), .Y(
        \SF2Project_MSS_0/MDDR_DQS_TMATCH_0_IN_PAD/YIN ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_15  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[20] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[27] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_29  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[5] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[12] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_11  (.A(
        VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[16] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_22  (.A(
        VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_SIZE_net[1] ), .IPC());
    sdf_IOPAD_BI \SF2Project_MSS_0/USB_ULPI_DATA_0_PAD/U_IOPAD  (.PAD(
        USB_ULPI_DATA[0]), .D(
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT )
        , .E(
        \SF2Project_MSS_0/MSS_ADLIB_INST_RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE )
        , .Y(\SF2Project_MSS_0/USB_ULPI_DATA_0_PAD_Y ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_9  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[7] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[14] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_23  (.A(
        VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_TRANS1_net ), .IPC());
    IO_DIFF \SF2Project_MSS_0/MDDR_CLK_PAD/U_ION  (.YIN(GND));
    sdf_IOPADN_BI \SF2Project_MSS_0/MDDR_DQS_1_PAD/U_IOPADN  (.PAD_P(
        MDDR_DQS_N[1]), .OIN_P(
        \SF2Project_MSS_0/DRAM_DQS_OUT_net_0[1] ), .EIN_P(
        \SF2Project_MSS_0/DRAM_DQS_OE_net_0[1] ), .N2POUT_P(
        \SF2Project_MSS_0/MDDR_DQS_1_PAD/U2_N2P ));
    sdf_IOPADP_TRI \SF2Project_MSS_0/MDDR_CLK_PAD/U_IOPADP  (.PAD_P(
        MDDR_CLK), .OIN_P(\SF2Project_MSS_0/MSS_ADLIB_INST_DRAM_CLK ), 
        .EIN_P(VCC));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_6  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[4] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[11] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_285  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[8] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[12] ), 
        .IPC());
    IOTRI_OB_EB \SF2Project_MSS_0/MDDR_RESET_N_PAD/U_IOOUT  (.D(VCC), 
        .E(VCC), .DOUT(), .EOUT(
        \SF2Project_MSS_0/MDDR_RESET_N_PAD/EOUT ));
    CFG1 #( .INIT(2'h2) )  \BLOCK_INTERFACE_I_MAC_MII_TXD[2]  (.A(
        \MAC_MII_TXD[2] ), .Y(MAC_MII_TXD[2]));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_254  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[2] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[14] )
        , .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_154  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI0_SS0_F2H_SCP_net ), .IPC()
        );
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_55  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[9] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[16] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_228  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[26] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[38] ), 
        .IPC(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[50] ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_214  (
        .A(GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_AWSIZE_HSIZE0_net[0] ), 
        .IPB(\SF2Project_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[2] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_114  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[6] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[3] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_108  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[0] ), .IPB(), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_51  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[5] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[12] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_238  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[36] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[48] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_222  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[6] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[18] ), 
        .IPC());
    sdf_IOPAD_TRI \SF2Project_MSS_0/MDDR_ADDR_10_PAD/U_IOPAD  (.PAD(
        MDDR_ADDR[10]), .D(\SF2Project_MSS_0/DRAM_ADDR_net_0[10] ), .E(
        \SF2Project_MSS_0/MDDR_ADDR_10_PAD/EOUT ));
    IOBI_IB_OB_EB \SF2Project_MSS_0/MDDR_DQ_13_PAD/U_IOBI  (.D(VCC), 
        .E(VCC), .YIN(\SF2Project_MSS_0/MDDR_DQ_13_PAD/YIN ), .DOUT(), 
        .EOUT(), .Y());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_232  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[30] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[42] ), 
        .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_142  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI1_CLK_IN_net ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_159  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI0_SS3_F2H_SCP_net ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI0_SS1_F2H_SCP_net ), .IPC()
        );
    IOBI_IB_OB_EB \SF2Project_MSS_0/USB_ULPI_DATA_1_PAD/U_IOBI  (.D(
        VCC), .E(VCC), .YIN(\SF2Project_MSS_0/USB_ULPI_DATA_1_PAD/YIN )
        , .DOUT(), .EOUT(), .Y());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_35  (.A(
        VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[18] ), .IPC());
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_119  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/FAB_RXERROR_net ), .IPC());
    IOTRI_OB_EB \SF2Project_MSS_0/MDDR_DQS_TMATCH_0_OUT_PAD/U_IOOUT  (
        .D(VCC), .E(VCC), .DOUT(), .EOUT(
        \SF2Project_MSS_0/MDDR_DQS_TMATCH_0_OUT_PAD/EOUT ));
    IOINFF_BYPASS \SF2Project_MSS_0/USB_ULPI_DATA_4_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/USB_ULPI_DATA_4_PAD_Y ), .Y(
        \SF2Project_MSS_0/USB_ULPI_DATA_4_PAD/YIN ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_31  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[7] ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[14] ), .IPC());
    IOINFF_BYPASS \SF2Project_MSS_0/USB_ULPI_DATA_1_PAD/U_IOINFF  (.A(
        \SF2Project_MSS_0/USB_ULPI_DATA_1_PAD_Y ), .Y(
        \SF2Project_MSS_0/USB_ULPI_DATA_1_PAD/YIN ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_279  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[2] ), 
        .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[6] ), 
        .IPC());
    sdf_IOPADP_BI \SF2Project_MSS_0/MDDR_DQS_0_PAD/U_IOPADP  (.PAD_P(
        MDDR_DQS[0]), .N2PIN_P(
        \SF2Project_MSS_0/MDDR_DQS_0_PAD/U2_N2P ), .OIN_P(
        \SF2Project_MSS_0/DRAM_DQS_OUT_net_0[0] ), .EIN_P(
        \SF2Project_MSS_0/DRAM_DQS_OE_net_0[0] ), .IOUT_P(
        \SF2Project_MSS_0/MDDR_DQS_0_PAD_Y ));
    IP_INTERFACE \SF2Project_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_150  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \SF2Project_MSS_0/MSS_ADLIB_INST/MGPIO2A_F2H_GPIN_net ), .IPB(
        \SF2Project_MSS_0/MSS_ADLIB_INST/SPI0_SDI_F2H_SCP_net ), .IPC()
        );
    GND GND_power_inst1 (.Y(GND_power_net1));
    VCC VCC_power_inst1 (.Y(VCC_power_net1));
    
endmodule
