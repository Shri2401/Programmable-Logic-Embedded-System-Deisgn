    Mac OS X            	   2   �                                           ATTR         �   _                  �   H  com.apple.macl      �     com.apple.quarantine  ���F�D೥m�#rb�                                                      q/0082;655f895b;Slack; 